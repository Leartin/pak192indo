BZh91AY&SYK��zB����������������������������������ӗ�����9�� �{U���V���t��[/o}�ύX�1��LZ��Y  UI���� W� ݀�Q*� �- J����A@�        '�>s�\��(�R��r��P�B4� 
=�� ����w��/;ˀ>�y�2�̱#��-|Ʈ�������������&v��ô��w������vP �.�u�"����Y%�a�L���ڴ�D�� 
J��3C �۾�n�@ ���I��ؔ��� ���D� E���>�m��q�Q�b�@���]u�Ar�u)�ZaQ�:�[��@ֆ������	HW���u���UT$Q�QG����� ��  ,w     s�V���$   	�0 �FCM4  FLL� & �� &LLI�ɦ ��b�D �  L�  &�	������F���鉁OS�M'��b��d��$�Sچ�hf��ڧ���O�3I�='�)�xS��<��jjyM�m44������&�4�B`����hi6G������i������C�P�=#ChF���5�5=�~�?T�{F��m&�)�z��O�=O(h��Dz�F�OT�"���z�OP�i���2�i��@i�h � 4   �          
JIQ�i=O&I�7�0����؀�&Ё�4@i�h�4=#�44hd z��Ѧ�@�d     "I� 	��&ɴ�hɦ�h x�M��ja2`�i�&4§�xM�ф�=5=2L��4jl�i���?����ښ��J�h�X� dD	��δ� L �-�LRF��y�Y���^�!�9��u�����2xpA(�}L]��}��Ƈ#,^�ts�sRd`̐�꺄���ZV7��*�%��*A�W��a�����^;`�ZJ�>ŌA�Y�Z=�z���I�W��*<��#��~��ܾa�k�bV4�N�J�b1Z5���0"J�ĩwJRbm^�yƩ�%�1�"9B�6hb��݉���&��	�Uz$�T+f��0���,KW�֩�;��\X����0�ֶ��+"�
��W��c��@�*�q��G�I���������m$��[�/�c�6�}E'�9J'vE)$�j�˛Y��ϩ@JP��G��w����'��c�iWyl��j҄��y�i���P�~
<�صw��3Q>%@���Ɣ�]�w���#�=��.�[���-�B��AX�:�mx���v�������}�L9U��>�����Tx�0�,��M�;�Y�&�% �����f��g�3[:�2�KTឝunm�;�k��d�9# ^<�o�IǱ�t���uW�8jbt?J�������[�CBֆ�֎нlB7>�{k�!!v�[t/Rj=�8��!����7=��!o|o(���-i�wVY��!tk�3uM�K�m�a� B�juV,T8��Bk嚸>ԉ��gC��}�����GW��������	&:��hdb<�d��d2ѯ�V�_� ��d�ƅg�����pq��b�X61��D�N��&�*
V	?@5Mi�sp�JVJ- � b,��2�CB �1�z5�p�)j��d�O!(�,���kiy�*��Yn�a��W��=��X0赱��� �{*�Ah�����
1���OTx
�П�R
�'w�㆝� ����I������||iv?(j��<I��<A{<��GS����9M$�h�-o*y]��g���������˧������k)��(�4�@�H�BPl|_
�(2Ө�\��X�˂���� �ޏ�?g�y+��7�n�@8����E��Bx��ڪъ�5sò�CA��/��U�iyg�&z�;��.�]s�����0�9E��c�{��\Id�\X��o�ӏ6�Fo��X��oY�i�7��[Ub����z��ܩ��1���UD�����SHڛ��;��B�{����<Z��,�=rD�E����AA��?਄ �g���v��`f�<_�V��5 ��&ɧ�/�}/�1��kv7����[���g
�M�7WY��K����Ϙ���ѫh��U�:L���m~rK����O���G�<y/�����5X��XjZ�h�V���G�"��r�
��F`bd48�J9�G6��ϫc����/<D���+6����=�L0�*�L���o{i���i)<r���.���ǹ��n�Ǐ�fzzh-Eb�7u�cدn]��:X���XZ�R�i��z���w�����\�Uw����餝��7�:�ч5�u��J�}�x1��a�����K*���L����~	�����O/�:�v�=[hO�B (�����#���:��ool�[f�)���'hvs��7�_B��z�}�����v{��K��L��O�2ְ;O��f�>���g��H|.�3���"��}��Ԭ������@ǒ�	~6��h��>I,n{�~ӵ�<���kg��[�oE��`���H� �jzl��M^�4��K빋;�_�sa�}>~-
?�)��pQsi��VܭN��6w���0*�\Z~�CC�sa�>����S�����fO���M>����v��|�s���njs#�7��l0���i\�-\~G��w�WZiپ�[�{��ڟ�v:b������'��]�l{#������2& �F������G�u��pz<���3��������C�0K������tl��X�,�2i��oZ�/��n���/�tӪdmP�M�������N����+�l�~_���G7{��ٙ6W�FS����-���W��k߷_MmS4���Zq���y�<��(BzZ��珞~�P�*kn���̺I�K���N��G?;����Y���������_Fƈ!��Ez�����i�x|��oysvo�_?�q,��*��X�2z��n�̔m�JE6a�{�"�qc,��:�4�����h����.�12��1*9S����;{;�H��uq]�z*��������j�<�T+��i|E�kd<]���K�o|�����A�ju<���J�^~�������\=��۾�/�Wz�d�����6�vpD��TxjL��)!���z�?C?c#-��+�Ǜ�	Χr�T�B;Y8<~���|*��s�A������M���T���u��1�B��g�����uw�����YQ�~[���K����44���aȦ�E]��z�ݽm�}܋�ٴ�{��mڥ��Lܹ�?�x���3htx[ی�}g�+5t�V�l[���`���6�f�O�8(y�1�CU3@	 �A�!6`]�b63�2X@I��Ʊչ:NF�������.�v^ǖ���z���
<9		�@����y�l�*�Hg�Kª14�
˥�h�ְQ����d1M�X� tp�XUT�<N[����<f�q-�r��4*e��^`���\���Ԏ�M=nr�5�[��B�zN%clh��׍b�b����k����q����
�$�$�����_��� "��r��Be�D���v�g��^�4�=�ej0�b�t6�N�V�$���v[�q{&��M�N2Jb:�&�����U��^Ds��M^6�?���U��!�W-SB-?zJ^_���x����T��?TXD[M��{i���b<�Q�����m�A8��"�%y������a�|��������&�I\�URCy����xh	��+	4)*Vn1^B�寧``���{}NjbJRP����Z�m0���dF:hA`�?��7��oqn�f�A�O�@�C�y/����M(e�E̑��"�$����y��:����C�W������� 0�stb�K645���b������{n4.���i&��ĘU���V�.����.B�a�/.�����$x}�]"Ap��H$poY]���ӂ���k�� � GEM����(&���������jT�q�K'�[o�a�hh8�W�V#eI�0��S��m`�Ǚځ��I��t�(��#��`0�BM&'oQ����ڨ
7�"J�_�p�N�#�dB�� ��ρ�)��1�{4���j�����a�g����y`�7�,�Ú���v���q�<�gd�2��۠�x�\�_�R��e�^�f��;�hs{���'�b��[0��_J��ّ|*2+L�7���_�nd�;�8�UU'��?�s��3.�X��W·�k�|Ȫ�X�䗪��}ZCL�Ā@{� �{<�i��U)��˿�����f1�M�>/�SW��DU�j�Q`��,�`lE)��̀P$wwF�����z�w�Gh�xu|=>$�5�ѝ��v:�_�������v��*c�xp����b��1Nj��w��×������#WU�i�R� ӱ�S� #���D�����Y.'=HO�7���X4!C.�o  �pߚy#@�v�'�9��J�M�^���5���̦rF��H��1�</$��c�x���������N߾�r��.�]%��^qXdy� ��DI= �r'����I�4���w���/G?i����,Rh��8�)���w���[y���T�PP�t�������������	�{����zO���,"S�����Z�+�.���JT���*�&�N�����*�sk0�r�0Џr����d�|M��A���w��|H@�Ld!$���
��0��|�txY7K�(7���H��nxv7��%h0��G���2<
O�Ѩ��17��'_�+9�������f��ۅ2^_ǕD�U��v�t��W6Mm
\MgH�;��Z�p�E&�����F��4�t�i�xpC�屣�H3�6^h,jg����=({�"��z{��8���e�'��Z�A^���]���ܪ���<��N~���uJL%� �������g���0?�J|�x�4���3�gy��i׃+�?�T&)/���^�N�*�� _��F���VdC���`�<�bOh�ػH�W&4�js�Y�_�
�8����^� ��F�"����
c��Q�~���^�( p0� 3xU�����		!Ikq����u� i���w�#]�3m�_~�ʧ	޻�v{X{�&鹔Z��$'C������M��௷f1�c��;y����.0�9�aL���jC�`V�,�R0L�����^� �k�y����@	�����퓉�����wW�;�D�P�����qv�_L���x��!{�����݄�wIu�q�]F�l�����C����&8����b�̃ �G[e���&� z5���
�y��-b��T�)t�7�5~^&����R�ë��5����������v�l�f�;��>����#��hm%��	���w�G�_(�4�J���3���7]q�H�	JK0M9g�����?����m��+ Xx��=�x�����s�,���a��_{5|WF-����z>!�+���O�r�$�7���mo{��t�2D�&K@=g��h��+̅�����/6uڦ�Ph:��8� �u�Ss2�e{,3�^��e�͗=�ɓ�X3ˡ�� /b��Š(x�
�Uqp݆���X��wiK�/�(��۴|gG����g����*Jܷi.��m�h� ���;����þ=���������|(W�}��Z��3`�Q�a��o��>�{�F*�7��!S7���ұb��h�`���Z��[S#7�M�W���� ���td��nex�����z��xq�T0U�lG���a����~T�yǁ�A�H���AAq���k��{M�'s3�&����:y`�BgИ����]�fF/�����&�%ᶈR]����8X7�.�u�<u5W1=*n�o�e�r^�s�i�A������'m"��Ǌ�޴KX�]�X�ޘ�Q�}�
]hTWw'^���Gck>;��K�R4&�0����}8��CEhU��m��@B��>'9����UCD)4���H!֩)�h��ƚ2��%[&�|wz������MeAN$T��@��-����}zw�k�K�3�w����z&J��Y��#����\ʔ�H��mid�tl�qi�7Є o�a&1c<�Js�j�f,7���~�d�HR9��c�mȭ��jLn^<�1�^KV���<FG �X�c��51���z	�ZM
JRHR� e2j�⭵{<1������>��b&D�|lA�[T��VU4�t���,9g�p�¶Kp�Nv�_	�M��"n�
-p4K,z���ߵ?D&���/���7"� P�}���8'�}��ny�_?rg���#�3�]k�e��^�I&�;1�Ja�ŧrIȕ!7�=��p/(g�~u����W��z5��r�Lڱir�|j^���5{iH�^���4���}��������ްS8�=c��{�^oyiA�!NZVfjR��7�9�`�Zu�m�n�
���m�rtG���Xr^̻��}�ƕ7��W�n�<.������^;{X4{���<2LG[����""@��~����>!T�Ϡ���	�(?��\����	��_\��(��������5좘-	\Ξ-����V���#r�G\�d���֬�e ��}A������(�{8���r]���̊Z�#Z��姹��LM,��iM-HӺj�i�hj��f��Qk#Z��tP��H�����oS�,������;��c���s�J/��U楤Ͳ���}`𛵥L7�?��2r"oGٱ��g�ʪŷcO��o+�z�����7�30#�/����ل�K� �I��J9��\�U��' ��m!��[P0�S�������R�c�u��+v٨��[�Z�㋜^u��/����/RLNI���86��8��2���{f^X̼mE	'z�gw��d�hJ@�%�c��y�J�9m��x=��s�ݜz#���5v�))X�OV��i�7����E<�q�,Ѽ3�Mbҽ�﩮Zh��>#��x%r���H0���#0i���ˑ�D�/k�Qr��n�[����Z��ǱE�Z|1�;[����\q��i5�����!�����z�k/.WP��1m���ܶ�4L��bG�ڪ�=���Q��E{�o���zJ���Y�x��&�z�UZم�a��ʐ`��y��f��`��<��f�n��pFitܵU���Ƌ������� ���\�\��݂��>1>S?�r�c#��kË��v�M���#Q��BF+�wt�&k8I����MǬL�Ij+�G"����g,���~��Q,��}��'Zy�H l�v�������=���B֑�e�-s�*|MJ�uŏn�X��:�#�nMq��6�Q�%���-�RI�R�i���e��]I��m�o�4��eP j��{�#���\e�TR�k�5�O��S	
�U�e�>Y�0��]��	ˉ���������n3��
��_�)G�sV�		A��LbB�\D~a��?0s�z�Ҕz��[�^����e|-�ӊ��jr�\G��p��v��5��qp��X����k�sf��&H��5O\\��2so�b���9=/�O+\��k~BY�V��l��������z�v�߰g�o�q���,v%o������~��@�y�vX�Lk"�M2U�Be3�/	Ӯ'��r��N�,$��4-�[(	ce5/lb/����Ӵ���)-�s;���[��x8�!��#��x�:��<^���x�V""��[G�ߙcTd�XX �$(�,�KhA&�D�/]p*\5�`��o�s�]]ʵ���mZa$�H��Z�VC-A�0�6���3�y�ϕ6�RM�]�%����$FO8��BLL��[W-Qx����Ydm��>bQ���Â�+nF)A�/K\����� ���`נ �9B	��bE�j�`�R� �
T
.��3'{�9n�14�C��(*��N�+\�D��1H��n	��1z��c*{�)h���mF����9�l�"��X�E;��2e<7��:D!��%Jz�C%'���Ou���ZU�N�e�r��m����6�x�6� `6�s�V.d-)��5��d��%%Z�&�	M�*�򍉡SLh<
�̓��"�#@O	>t�)J�I�8�I���s%����@�)SΙ�����=Fl�4��rփ�(D:	-�ҡoky�9�s�q���Ƣ�6����4it��;���M[S�y�� =�p��h5���ɖ�������v���8����u���q/��;T�%d�|֥�=tӂ�+b��խ)�$55�t���
3Ὦ6ɷω�n"�;����kgek9��9dp�[�E�2��g#�#��֧����yW��\68F����L�
��Q��1��
SaC+A�RzMd���=h�\��sFw*0I�d��X�scrk��:�O��/��ޮ���{ލ𬗫B�x���x3k��/O"�w9}s7��k<q������7��ư{�޻g�]q�����k[zŖtM9�u����;d뇓���v���<��z�̃b]:�6Lgjc��=�9���,R��EnHrJR�5ϥ/rԣ�iq��C���0�[Z��-ȐM�i�^��t�m���"��hK�	س7�Km�W'�<+R!:�Pr�D���f>
�	x�eRo�OD�������M,m,�Q�Rh�S��oS��c��&2U35�l�ILP�S%(�=MK��)"��L���"!��"3@�����jb��,m)�3O �����S5�{$J�ƺ�Гc���(����[ޥ�_:օJQ� ��)1nZ�y����1[�%����u{:ļ�Wׁ��[�^��H��h4�	JP�6�Ǜ��9͞x:����Sq�U�1��'*�b��`���]�����g6]�p�O/b8���{j��c�>|33yw��w�����%!�w�5J��1�J{` �����?��i�5��6}����ܿ0~<tò�� ��^#$���9DLE/4�����u�����f6E����n*��/����6��7�Q�e�]W|-o��=���O�>�	���Z����3g��m<��Q�䂙������X.j���m��K� �䵃��,��UTT�9L"���Z�5���]���q!.%�SO����Ѐ����kH�&˗��%)F�T����W�����c;�����X׷���O�?�}��<QFI�!Y\\j�z�2�1�x���D;X<ڻũN������w�������Tpn�k�o_���$�86���Α_=�y��5;�8o%��h[��N8�+rS�Ŷmv~,8�K���t4�:��͍� �C1*$ >sl~�	��952����N��O^{&QvH��Ē�0��BF�5T%�"0,Mj��3JJE!E��"�$�B�&��N֯*W�m�ňIR���\�	�J�*��&Xz7�k��=~�O���!�2���i-4Tp�f\`�����.a�g&a��&�ca4�a�C�ЀoAr,�R�P5�%y���8��2 �(�����F�-�  k�����MO��?��뤟e�{���R0�%��
��XŬ�=�\0�E�BB^9��M+De�w6|��	;�zI�f��B�{��ĩ�&�������(v�����D��t�TĨ�QE`�@�8�p����q�������5.����0������	s����}��w�j���²h!��@�N�B��V�4�!T�s�6���6OK��,�Yt�0Y5ϋF�˞L���y�_w��
���a�(�kD�b%�W$/p�EEwi��n���� $�u)�� @^V:�crwZF�n���+�񟻛�B�{V�' M�Ѻ7�naU����d�#��9�Nu�g��(��V����$�f�CA�}�nׅ�?��oOd�OSQ�z�UoU'�v���p.�DD�5J����B�v`?���bD��#@#n0fI������m�a��q�h�^��	����H$ohf��	o��l��?�b�ܚ��p����3��,� 5��9�N�T30�����60o�{
]�y��j�����C.�7�\|N�^�v�[�6^�3߳/\������ʹ0mIءw�T9.eu��q?��3C��U/h'�}~}s%�!	M�5d�O�R���*�>�X�Z��,��&����ܞ>�R��_��*'��Ta���c,��"� ��dt=ut��?�n�_R�����٪K<�{��x��u'g/����s�7P���}^ۤ�>�&��vPF#�0@ �����E�DB�u�˄)s�3)���/�\���C�].�z�[TӤ���P�9�ҙŸ$�ɛ|�k�2��i�31�Z��y��t��^6j:�ifg<��^:��$k�=�`��zr�S����w�~�!���9f�O��]�|�V��� �`�D��ax�L|�����z,�a c�~�"�T+����L��tt�L�=��ij�v#��"� $�"R?I(�uГ@�Iv�=�D� "�� R��T�"Ҕ��1 5�?ߪXwM�&�ẇ�w����ԳziӃ׃�Mi�_�4�(���*cSU������j�x���
�����5����zEy�>�<GW���	עrU�^$k���Vש�W*����~�u��*�.�I����O;�7�&��̵?>�������4]����:U}��gbםjz��Y�uO{��,{?��|�SG���B.�L�2Ԛ� >��/7Pn['�a�h<����?Q̔UC�aE�u������8k�?��Z���y3#h�}���KŞ�g��@X����t�����3O��J(�~V�ԣ�������a��R`kB������[H	��W��'�$�QA��Y�ҶϾ���@���uC�.�y04��9nw��-�p�8:��8�4E��1�J5 ��nؚȌ��|���Dц��8.�lXÌS@�hC�J��䲹U�/�e�w����U�&��A2��D���ڻ��b�7	��%�$��d� f��E��?U�k5Cf��
<��?�uI`J|�;��K}�s�$�.�~�������Boߛ�E��@�ȉ�4eLS��3#�PB�&̄!���)F�u���&�?�r(�b,A$����T���v86x�6IzJq��Û��;?���5�3��1���xJ<_�B��@��@��h�&���J	8�@�m7�t�16�:q�J��H@�BҤ�ޚ҉yN����k��%1	T $��UV�@MՂt�Č���N���7����:�o<����7%�]ztb�v7e�1z;��	+�^��h�V1HĪ	�*#4ܤ(Л�T�c�e���r�5��yrkv�f�OK�����*eSBE��L�Up���it�ˑۛ5zoM۷z]io4ɂ��D(-T�#i�I��$J��ۉR�jQ)�D:��T�j
H�rAB0��n㑹LRH�T�Z"I&�b�lE�A�AU@Q�ƨ�D�ܒKC��I$%68\b����Hʻ"�rJ�GU�jZ��%�E#�J*1��Z��SBAm����F8$))&�c#TIE�A*CM�mԍE �#N5���&��F1JCt$F��!�m&(�"j��81� یq������D����!6��IH�!6�R6�(1ۦG�v��"ۊ�5Uj�Tm�����$�#dPm�7!"�������M�T�AZM�b��h�$�j�(�BU��ҩ�����ISڏǚs�0��]�]71�];��*Zi]�9 �!�J�R9	LqFB	��A����H.�D�X��ն+CJ�Ub��(ڒ�$�N5BM9$QmƘ���I$�#L��8�T��M����rF��nF�J�!��]�cZ�ɵ[��4cI��e�v��"�\�E!��t�wTX��We%��]A����ו�f�S=�$5a HF�\�^��l=b�n�B��̵Ii@�ku5�׵�]�:uλ'1����m����],q�jcK~��̬њ�i$h�4��3f����"@�T�h�M�[	X�$��Km�gʧU�;�%��U���
�6E8؊z�	�<�y��ou�1�����A5 �z���-UG�����z�_�#�1D	O7���*^���b�4F(��+��4���c����j�A5 #��P���Y�=/��q�*m /��M�ֻ}v�꼄�`�mP5����U�2 ����6�k�����O}�E;�AB�AD55��&]
]�V뷺55���)sAAdC��]e���"��BD(�ϑԣ��*䲩^���/S��v�H��E��(M�P�	4"�&���<���0A���.`�b�4S�5*�-��sr=f�*���TB�M.60ԭ��d�1��ܬ=q��I����M�gK������8y��ܳ�MVy��u���2t��W\��V���R��Q0�ĿU�(vՕ9i��˕��#����/���@����_��0'���\�<�E5��������m��Ǐ��J��M*�[���QGh����8j-��k�չ���),��ٺ��=�V�u*��&:���t����" [�a>�V�[����`d@?�[Y<e��:��幌��Z�v4z��֕w����-q��Z��;
��g����G�L�N�f�T�jn�z:��	3+|���->WLe�#u�L�w��&�����C|d����.�9ב�u���M_���DU��ܲ���4�	��{�YZ�CM6-���O�7����UwH��Z�1�����ӑ�-�e(/"-'��Ńu��'�&�@ V�%D�&4�DT���i��4W�}���_l�D@�����g�5R�Y�Ԑ@"�+���� v���h
ku�G������犖�$��!! ��f�����Ͳ��:|W���:S`dٖv�3L����i��B 7�.�mu2��i��o�,��s���ի��eu�z���l5�FA$"'�嵎i��]���Q3�x�	�����s_��_N�p28߉�^�� ̀3&D ΢R�\���j�iݓ��A�nqc�Y��e���e�fZ�[(��LغZV)s�Ũ�ۻ3�D�-g$Թ��/?M�Tϥ��댚
+F���]��&���hB�,��R@�F@� �(�h[�X�tT�u��B@	�$d7Q�E��zepgө�\H4�B�y����o33j#?N���Nei�6 �#3?�l��Qc^@�0���끿F%��N�x�ͽ�B�Q� @e1�9L�Ȁ^A]R�w� 6�[|�L̈�g�W�[���gL�8l�����_H�!�����c��ЙK�7�	��?ECGu�S�
g0 g��[�P�Q�uok|jDd@b�T�~�筵�� ̀ÏqU;p�!LR` M�ɧB�2&�<��s��� ff�@9s;ӭٳW9�>�ڤa�+M�$Y�A?�ٌ2:�>�>j�
Hin}�EV��Ҽ�:�L$	^��٫U��30YZ|zѪ��-	'$�9�߸�Ȧ�w\���7�(]l,�.�������
���e���d
[��r�+3����@bv��+���]|9ڛ;Y����^� �ᦜ�3&�!Fr5��O�db�h�ҫ^ 喧�'���h�� ӷ�ū����۬�:��j�6���#Uδ,_ǳS�S���DKy[��zx0X�������(�6b����B��x�g.:�[%i�����ݾ�wnBbTj�nXgW+�|Ĕ��f�>T:�>�w5o�43N��fyȀ��[�p�����K���O>�ȳ ܟ��	���0�0aU�ҵ\
ʈ�"� f����&��u,��D1�g����F�dڇ���*�f��t��*�t�vN� ՠ�e٢��rQ�h,���$�L��o͡�
����1'�V�A�#O~��N��خ�[�k8d���dG�%\�&���N�(�Ҝ�� " L�Ne��@�(�o � �"�E{�h�� �M�6p����d6�eT�Q  ����Y�z�?J�|vD��w�x]^�˩�{��,����m�͟-�9K�柘��=��z��ְ씑�*i^o����b��X�lFVMD��}8�G�tF�T9�~�L��u�A��Cs����(�|UspiT'�J��̓"�7����mv�h��:U�P�k�;G#]��Epp3Nu�{_�>�ħ2/Ypjxs�\!�-�4����ߏ`��N�9+g#r�3B}�/U�NF÷my��8��!ߌڏ���\�82(4�Gr{\������<�SO;,AL��(�t�.1dc�� J����S��Д�d�6ݸ�	�5r˺����Sṋ��U�1'�Z�vl8š�y^�����1m�c3�.zx,E��S�.�q9��ե�� )������y1�gI�/�F�2�=���7\�r#7
d��7R�:��dr���˂9z�l�h�@{n�"&s�
��3C�rc;CjϞ���vƪ��D"�C�-~L�lҞ;g��$��lڧ=(жW2�۵}%�6�W�0U��gi�6��ŃCa�"3�vR��͙Sc���$u�G$fЄ�8����8V ��\�ѹ�xoK��v#��=<�VEw��Lg���6`�<O	���2�o�����t�=Q@;�u�U9�[\z���tI�~���O_4d1����Ȼc{8���t��ܥ81k4ѣ��4�v���f� ]��+�<'і0X:�I��S����ګNå�>��:@�\<}�FV;k�x��A �̇) M�"L�t�.HE�����;��e�jSC�Wx2͙'S6���%TȘ�����Ѹz��9
k|Q�2�<�,��S����/�}r_[�L0!�]N�!Z��ÒS��<�8`��F�#��g���sk\�>2�\:(�b�� �A��P��IX���#�磮:tf��C��O�S�������ֆ�Gk�Q��"E�K;�4� 1��տY�S���S[k����c����Y�u�@r㮣���9�
���S�ih��(6��;gP{Zn[�3���a
����}��DH�#v���UXU�KXj�O���u�-$s⃳t3� �ۺ��L�цm@,����%��[> �a�5�4�ϧ���U6�-�W��G�u'3i��t���DME��� Æ�E6�)��.�Td:�hb�&��f�6�]�ȼ�`x�E�βo�gW:�m�*�@j(�*Ƚ^�+M� :C]Z�&���Y���0����v2��ֆ��� d�p��k{�n�8w�����/���5��Θ��D��ڣ]���U��x�º�Q�O&�{�ձ`Yi�h	�Z�M~&;k���Hor�Mg�|틔�I+BƂ�����xEwPɼ�z�EH�M*܍)uʣV�p���s�.�#ڔ6�M�S�}�kb������`�F�a6g��<>7Li(��������8��`�f�^�v�|l���<�{4ld�ڳJS�&���7ve�$6�w��M�my��ٹ�Q�\'�l��_�fL�΅f�㩝tYB�*�/����E�r�}rCk{��6�QfJ�YP�DC��:�^('H��t�K?2W_�ء�M�5N����ӮA��)���Vֆ�(e�����k��:=�>�E���r1Ƣ)�[�0:�\�f\r�Bm��"~4����3"�U�Xں�eݚ�3{K�qǫ廲�F�)΅�G?J�jet����ۯ��^�ޖz&̉�T�T7��I�A�.>����+{X�W�l��)��u�(��gm�u'92�cUlD!l��kQG���݌����"��a����*9�1�����	��dC���3�j��-Z�Y�[��ꑓV�.�a��'F o�Uz����J,�sd�{����'o��8)C�F
(�i�bqHE��D�s3=Yv��������*����GqR� ���|1c�r�J�,�Y*Ҿ��:���Oaa}��ȡD��C�%�=�o����)�4��w��a�G���	�m췑����޴0S�����Bf�`�2��H��٪�m�ꧏ[^Z!M�
��Zy�a��M���l��\TP  �" D3m4�[�6��+��~�q}Ѽ�_w����_���k��{�2l��"� Q;�"+��Qr��[�p7�V�'�n����5-��Ƶ>39[+J{]�4U��B����	d�C��M��^M���|F��u9sC��mX���p�iV]�٤�L�z=�Uq;r�
*b�=�t�E��
ɚv����T��CB-��U0V����[�j�_E�����T5 ��]X�!*k��@!�M�U�D��nk�yur<x��nc����:�1<�y��k�4Q���b.��x������%q#\7�t^5wv�㻭���Kx���+�vȍ�j "qDP�(Ҫ���}q�O<���v�^75�oTmS��U촐����.h��=e�eU{�(�<|v��W2�nj��E֖�m��*��ᙅ
zYUG����J��Kjl��|.���M���W�4V�劝�dsD[�m�\���s;��6-J��F�r���]���.���ljH�,f-��]�Is���w;��$�77/<�Er�u�#lU�-�Q���#N�湮k�8�F�*��*�F�m�`�;�dw[��5\�d��W-$b�w�z��?�����\���s\�R�Ǫ�~7�_�	~��El��*4�kPq&��	ڨD����zf
�om����i[=���X-"���4�#LpY6G�z�/X�kR%5�apq�N/�0�SU�(z|mB�hUnFn�i$'.Ȓ" �sr
E'S�щ�[�RW�.+8˶-BbD]-.w�=��q�:gM�k��g����1����+X���"I����Ȍo"]@�c���/U��u�M�(QS��!���C���	�_E�^ӤI�����h�?ŕ�Cު���'��z��^�"��m#`}������m��n �������=װ�c�f�0���b�^������W�%Q{�^26��/�ʩ�O`2�q���������P^���A�U;��􊟊
)�����GR";�����{_�癨�ǣ�M>kP��**<]ܯ�fԯ��}n��q;�Q���'F	�������P��?�G����](�H�s篰����a��[&�"'��{�o	4,��Ź���|^�ܮ�'���t���A���_�`2�&Z:X��'/\LO!t�zCm��6~��mƄ�� 4!�"�kB�B'��଑>]!�
o}��7�C���wl����W/=����DON��_c�|_p���CA*x����Hx~�G��<{ ?ZF�F:��q�h�^������C���s~�qp(�9v�ӡ��M�%Hrg�~׹���`�x�4�� |x��_%(��Z�)����30x7�]�"&�'|�2J<� ��zsV�HFB[����|�v��k#�u����{-��bd!z �2!x�t����3���3Q���(�?;�D%��c��:$MB�d �ꆨkd���>ə�U�KL��yz�~�U��3|E�l�$<�e`7;���(����/e�m6=�x~��N4��p�%���n��4�`%#��V��
1�H	2#0����|7�ۏ<�m���Oޮ�U� �D��� �J�zA��=9��`,��@"�"��E=2l������r���8z�Ʒ�d#9�<ܞ
���pt���C��M�I� ��YҘǴ��+s\�'�HVD�oK�� w2B$$N�q��"{a|�lF����C����v;��ըt;ٜ��]�Y`�2�~y������!y�Ǵ��ؼ�X+�έ&Ub!�(v�6n�m�~#���A;��w���|'����}�c#v'%�WMj	��y�r�&��M��e�%�z�)ML[o�kC����K��W�g<K��i�4�'Inb�풋X]���3Ga�����n�6�Ivβ�H��`����(�o@ Zf�v������ч�q�����Ow��J��q6�#	}& ���|p���p�	�X��Q���Xw���������w�tX#�û�i�����g������27$)�A�C���REӁ�E<V������a��09Hps�r;����מ���y�'����o�<Q���p��spu�`)�<@9.��z�Yxs�yP&���� za��������G�C�C����A������Fm"����� KE;��i4���T	�6�\j@��</X���O!�nC��s���'�M�w�H��;p;�=h��5��������k ^D`ea���>a��o�˺a�4����2�h�@�f��g�ǣ��� b�E���E�?��ݧ�$�`!�G����G���M|�	�J�2D��1'h��D������4=���
=wk�.�C�� @�__��c���I1E��6���eo�����8 @j��r��������Ki�y�σ�nK�LE��y����'���c�J������v Ay�z��Q<����ѣ<;�#t�؇c���g�;ze�Ԇ�>��.%�^
B�[��UP�˥��8�b �>�rP:�L!�����7�8yzG�϶{N���D��𽴇Cګ��ԯ�(��K�#�&��0�y<J�8N�k�z�������%*^q�TM{�X �{�����S����I�Ǵ�~2�|٣��ww��Jj�\�h�VH�ϖ�\���Q �O��x��\�蠿R7�x�
�zՒkst;8�c����o��e�z+�:�}��(55iC�zZ�<��`1I��x���^�G�B�u��v���zi�p���x��r��^���;qW�Խ���ʇ�_�ݦ'�Q�z��=U�8ꇔ���TvPvq�9:|l@�\jP�1M~k�Z�����\k��x7+����8l�r � >5����c�ۓ�4tM(��Կ ��pB�8BT���Z��9�" �͒GV���$�d�R����V+� ��N���z���K��k��o�k"zؾ?w���}�UMn��pz���nP�@��@7�/-ю{$����u�c�0>`<�l1VF��!�g�-�t�׆��X+��C���� C]�Hƅ���^Z��K�A��OI��b�C��^����e����Ň�Pl�m-�D�e���<�b����Q��y;iAwp�q�I$1��І�+a�z�1@X����Ä�>�C��h��ge��C�q����|���Ҟn)��j��?�����op6�5�y��;��ҧS���$T�hkR���=���"��b��A3�� =�JG�A���}��m,������`��#�wр�Q�(�`1EOG�Ѧ����L 7@sE�V��M����{��y�˔����T��U!��zx(p#��z����!��]u��<U����v�#�ϧ3�A�<{�]B6��:؝��zXq�s���~Z��'��? �$���r���ob��%��m���7Q8ؖ����p:���
R\a��:H�*{F�����y�Z��+�l�B"j�G���+c�q'!e�!��QM�N��P�Ds�4*�79K+td%1A8��������y؞`<�h��zo�I����m��8�_p�DZ�<��>��I4=�����4 Z��ty�v��}M$H+�p7ކ�M8&x�
7S�*ա�x[+��G��(W���G��>|�D�S��5�CV,T//��x�3��'�!'���&����{�Ӗ��_�V�������炘��۬�l�؆۷�CpM���' �p�
wW_`I���9Z1�6'W���b�
���O{���n>-7��T���� �F�!
��m��r�@n�{}�Y� ��Q�s���@t�mZ˧}���
��_A�ڊ�*&�i$X�IҒ���
��h�Xն-�jWИ��')�6��[KiE�������[ؓj�cj�e4�xi&�ڦ�-�m��[*�	��Cb6��T9�F�l(�b�B��`��m)l��T�J[!�R�H�T�QF�#븃��	J7w�S��'�n*�Sۅو���?�'����˼���{K�8��z.��>�ߥ�}����j�PAF���K�|��,�t�
,	(�kܵ�6'��ޛj�k�ذߖ0�x��2������~N/��g��AZ�r�8��	g��7���K��t��z����2t6I�1�0�w�}?ʭ-F��O��I/�v=�,V��
ЅV-5S`ܬ�I$k�$l�.P��L�5��<�s��� p���	�C��|ߓ�U����O
?��/�O��������4^�6ʋ���~�7H���tXjw<Ug��ڥѷ�]\߃��y�~�G�|����G��]74p"n�%@�dBӪ�b�j�Xֱ���ދƱ���g3��"���R�����M2O��q�
[ �p����H~�m�Z/�v΄q9Rn<j��/5�������8���*���nR�X�"U5��k=O�[�����/R�ɧ�҄��L�2Գh�(����9����Il�Dﭓ��u�u�8��Jt-���%�ԁ].}[?u9i7�"�]�4�z��^q]K�ҟ������:�g����i<I������ؤ��_��m������̉��8�Ѹ�q�<p����#L�ŉp��yO�	󈲘����S��jl[��@�h��~�<-n�d ���ǒ��.�{8���!�1j0���%���e�Y�b����m����قH��<*�6玩*I+ekon��q�S�S}��*T��J��Ush
Pʓ<W���I�ܝb�O�j�#4l���fc/���dL@��F,TF�$uB6K6:�w�_%�ڪ�W2��3 �k����f�Yd��,m��%>����sf٭�ߓ�=w��\7&1�M��1�m��'��c��lb�-��Z�W��ʳ����襾0ƒ��tg<��\�$�ZmPGxĦ����p�6�mӇ̚�e2�l����q�f�Q(�j������]���ѢP��)�E�M�WM0�Jkz��g9^I���O�۶w)�0}�OUp�U7
��r���Ub�19�O��#�@�9�n��տ����������L2[�1�&��c���Ok���y]_ˁ�~!�c���П�ȱ�i6sK��oR^���?ޯ�m~܏�IOz�e:���������a*&�t��~����a:vϞ�*�ox�,݇O��+}��.y�k���~�o�eې�F N�f:�>�͍��,;X_�;����mN�S�u�� ��/��9�Ȱp�neG7��]fӯ���������O-W�\Z�~z��-�u���3�5�?K�u��mkW�k���z�_k�����w7�ّ���� �N5}�w�1Ǽ��j֫�&^���`�렯�E��)��̕-�&�3J����&�M���
���Uɭ�a0Yc[j5����ن$����*c��m�e�D%��AD��l�4�YV(-��V�̣��A�Ƃ�<�D*����J�Kh� ��� a�6K�2c���|� 3�礢Ȧ�рI !�=������u)r�� �U=��:�4.lZ��D@!S�{�]�ʀ�󐼋������O���xA�*���YOW����[̛U}�P�Լ�WܗC�^�"~?�)S�u���������΋�bX���1o��,���y;�f� 5��XS�(Ĭy���u�����������H�h	�b	� �J��*[llJsI�k�U��̒[��O$P��G�Y[x��+��omu��#H�g��&�� ���&<�� *#�%jdE58�/f?_���.v�+C���ێf�� �^"�Y���I�@��v��]���cK��JfH�~�����PjҒ<g���u��u��z� 6�������X�^�V3(�?�hߥ�G�v�9]8P�te� Q�!.!�� .�?�\p���X���5_���tR ��:�8FBL�M�̀���I��"� !�-�@�4"o- a� �� [�/�w=.	��jZ�:7�<g���?G%���K�~���p��Q:�.��`g�~6�g1�l�qJ��?$
6��'!:�{yo�F��=��+����.�ݻ�8�\��%)��|P���M?4	߻��e��H��	�[C��&���&S�H���B@ ��P`�{Fi�6U� `�/�$aۙ <���T*��\V�U����� �g�_�E��#|>U�w�F�1xjҀ�c��[	"Fp�\��<�ކ~��jy�qvSBo����۞�{��M�S���O��{ty�^�j<�k�'���O�w��`|�	�5L�/#,b8��/��`�(٘�?���'�˫������؄�
C��� &���㩳�[~\�� ��
2�?�w[��Aiم%�2E;�§�\������l����)�[�4 �I\�lCVpx��H&ڱ�Wh
Q�se�T ��	�����?Bbx>"�2"!6����uM�e
=@{�ڙ�������	5�*B�� ��M��,�?�J&���a�t	�E��`H.0)]���C��I١��իq�QN0`5Ȓh`�Jye�H�39���=+�A$����۔*���Nβ���=�r<Md�L�d.'E�X��ꡡ�[Z����5�=�+\RQ6��gq�̱�s��ղ�]k��tw�B�G�	���[,v9��=w��ء#ـ�����+�u���x��-v�sd9��@7����x�6h�"�������/����F�^R��t�&���+��?��z?�������.I�$�[�E��ԙ�FI�dh�1^�ݯh�URMVj�gLm��ۍ��墽�5��7m=T���~�~��E������@���q\5�ғ���-�u���g�a�Y���:����'s}�ICx%�)H�cT|3In�W4�M8��:"ײOO	�.�,�BFo����P?��~�>�j߶���}�a�s����p1��K�;���Z��[hjd�K̀��U��3_��ߣ<�~v��n;c˽�gKC�������N�NN7"cJ�����j����O,0��"_)�v��A��b`6��&��~�\`���x��س��Ǔu�LU;Lum�������mpv{u���лhm>E��7��m���Мq�C��R�D-�Z�i˶�QI�F���6�R�D�&�k�Z���h��EPc��p�(ѭ�e�ڻ`lf��m��m��$ly�" `a���:����+�w�T������4��Y[�m�����y̤�߁�x������o�����$���$�>Uv��v{��ɳ����� �k'ͥ��OGa�����l��s��oBh�5����]�L��=�L�3.���,��SØ��6x�zH�jh������n���~���{���t�z�5���ڿ�ݬ���N޼����csx ��D�FEW�|����l�l�o�����e�����ͳPO=-����e������D�Pqb������d�a]i+��=?)#�S�O�sl��ȡ����;�&���u,ʃ�OJD���ǌ��؟Tՠ�=%	������m6.n�����v���e�)5&=���KF���J¦�{�W�w7�&ʗio*��LXT0��|��0���q�Oŗ�bW15 ��@tb���)�(Q����!���Ϲ��BTy�ζ�>G�+��E�`_�]]�NǛ���4��~�����{������#����	 ���n�\=����g�K��e��4Q��wC?\a�=�r�=�u8�;s����� k������+g�F����a�J� ��r��-O
f�kCR����KU	�I�_��iG���|o�mԩ���L������;�������_�>���)�>��Z!9] ��;\,L���Ҁ���_ڽ�{�u��y���{�F�l�]�B�����M��g?'�y��`�M�������z���]?�|�'�Ű��ܜ�}�;(����}��D�w���̝����g�c�."{���M���B?B82�� J�Q��P(���M��O����԰'K������T���=���f_�;�{�nv{��6�����dm�=�O,]sO�����cm���h,�ɱs�o<X�O��7a��/d�)t��'��/��p:s Ed���括��7~����ٜ�}W�;a~�a���Y�@b�핊�-�4��wuͷ�U��ڀ��\�a��k]�M�Z�)V�h�Z5������I��5�E�.�dֿ-����ݻ�(�1� H�v�'���s(�B! ���T�I<���w�s�W������!���O�{��h;��d/�cy�h�{:�o7^�}��1 d[�ii~�>��pv��_�d�x푝�C���l����+޳���f3�kn�R��� N�����݋��{f#_�<���S?1q����mkl�M)e,�|d�$�@�N]tj�kZsJ�U�R拙J����\�mssU�̩mUm��2�V�eKeCk��&ԗ����y�[�FRv�քu����N�/$�s;e=��>�΅ْ��&E�����1�kJ�i	�Ճ3�(�HR�>�F�}��T����Bq����L)g��㻍"t+����0�"W���b Ϛ��ȯQ���{�K?޿�m�5Ry����=�! $�M4��RH�<���%�����y!�{~�CULڣ�R.����|�G�k�h )ݶ������-�眧߰����6?��F��j*�����ߐ��á�����<���O���s"4H�Aܮ)t��ыs���:lv6
�f��j��ψ|̻P�,�ۜ����7��߇�yFx�,v^�s_�D�V�:�T�KMfZ�s�̹�2�8�mt����:�Ѻ��6M��m���&ԒX�(��T[EQ��ԓ34`�m��/6�I�jﮜ�~S6�ڶ��̹�*T�P�R�G����o�������l�{��dU�-����T]%�[H�ʤ����W�^�9�7B����T#��o�7#{�����������z��e����^4���d:d�J� $J��:BFD�! ��͂�p0�E���49�S�]�T�|T䅨�����!#%UO�6��oD{����4���2H�}��	�WLa�@����kZ�$�M$�*J�̂��E+���u?��b�d�ot+*.-��m����)Z�6�F��r�]v�?��T=/�������ͧ����?��?E.�3�oy�c���d� ��3�l����`������k�2�2[k���2�^D��Oe��� b��u{w6o�QNV�BF�`�Ζ�4m�楩6��Қ��)����9I�T���Uh�h��i��F �D%U�Ո+YdI�REc�t�������k��?^���_7��c���]��������O�������o��k4NO:Gg1��Uo���%�B$R~c{���_�f;��..p!:�+��B�xNs�A~�ΘeLYF������?e�p��~/]�+Ĕ�z�Lm�l�x�v+Z�ʉ1#A�2�ro�՗��Ɵ�]Y:%��V��݌_G;h�Qo>v�>"|L���y�P�_�ǃ/������y�e�3_/#+1#*D  d%� �������)�ؚF�3F0TF�z*���Y6��m��Tn��AIDSE�L���V�j�f�a��x�}�-7�!���=0P7�<W�O�����O�߾�Z�.ju�{*�q\��M7��G��J�:�����q �X��,@?��VTt����ﱞ&u��x{�W[��BHJ������{';����������w~疬��OX^���+0�BZ��_�a��}W){������3ߟr����.=��s�Ҁo��1:FD-�6ɻ�"�6aj���ۚ"ʍ�h��W�7�蝼mEh�d�DV�m��r�Ll�9۬v�%̻j�a��*� @Tbc��W�C�'�_�����\��o���A��Z�g�?��v<��}�c��c �,��Y	0��J{1Ͽ��X�SH$��J�_���F72� (a�ԈH��^ɕH0$d��@�����q��/
�d�f� I�[�����UW=��'~�ɽ�w?Ǥ�\�}*}�����v޲�l>Ή�<ʛ�F�e{u��YZGX�"�F@�@ȁ���Mcņ��~��جQ���m���o���3 rb���� ���'5D��
���g�ľyz���}[��6+���sy*2 �`��⎏D��q��D��=��QlA;�S0�1!d�,���L�וW����O����T8�ȁ#�*���V� *�%��5�/ ��,CJ�$j	�
����Ҵ��4# fZ�0f��>g-��_	����k��:���8j=?6�.ﴍ���~D6{���T�ܲ��]|y" `�0��eE&�|km��(����Ȉ� ��q��X�r:�l�l�F��7RtA�g-��&��֘ڶ���b�9�Ѣ����PƦ���K[H(ٶ�)�h�5��0֑�8R�ܵ9��Qk��;��Uͫ���E͋t�&Ѻ먢�Z�ʦ��6��sI��bM\��m�r��wU��s���q�\���:T�4�%�r�b��m�n�ڊ�p�&�m�rܬlmr�m&�lk�-��h��[���j��rܰk�r���j�؎S��m�.\�ElY6Ƌssk�-\+�s[sl[sn[�sm��˛r�ʮlEI�cn[&�N��,X�lZ65A��Kd��QPEF�&DDdD����|�{/x�V�����:AD!��?�����Ū��O平���<ѻӆ��I��'�-A7����		$�I��Y��ƚXY*����)�4�8J^�'~���2?�3&�vqԽj3����Kd����mo�����0K��\��X��V,Z�]�J��j#kλ[IbFf���ʚ�Vk�rk�Pts���X��@��"4JU���}N���؛K�i6�cũϷ8�٪��J|Zĝڃ��UԨ��Ԋ�������O
�!f��X&�1�[U�KUb�L6!}@��
<����krytК�A�ϕ���".�vIH��ޝ���9�߯��=�#37�s��=�_F�
��A0`+I� �0ff@��(#����ʕY��f���|q�z�����w�v���s�m���d����!��7ԋQU�H�^ :�e�-�jd�����X�tP��E���
/SM�+��>�dLBf��$� $�n5+�3�K���!p�;��K{�����Q��x�������c1]۾������B!o2 ̌��� ������T��5܋�rݯ�� fF`��FC����Z��Yf��*VE�:��k��5�3��]���H0h�@�����ŗ��DU��u>�]h�B���JX12`�y��o�$!Y*F�pBI �1�պ�/q�4���-��+��;g����_��K?-��aU���`�7xhם��@.2� f@ ��! �0F a����:���BV\����m���k7���{������zAWr��w�^K��
A� ���^G���Tt�TpP_�L30Dcs)���w�y���dr��7��9�y�@ɦ�3���O�#����m����xd/y#��m�	V�{-\]��������/9>���W�!.�����A D`���!�q���}�l����W��>��M�y�k�j�>��ڬөb��k�'�>�XY n*��(*��?�dJ��+���p�(|?C������E���#�4�2h�Ҫ-=ϋǻ��������
cE1��5�d����'=x����No����\~�G��!S��m��Ih�f2 �� $ 2`���]wI���������B<�u_���m����t��6��G �բ��&��mGnʯ�EU�V-E�)�h�F�MR+I�Ɉ;r����9$�&�5"��_�j�9�K� �ֆ�c�LQ����_�p����J�RP�K�7e��W�k����W��~�k��k���sY���c)������iK��A�� !�Q+����_G�������6�Z�$x���:�<��|�e������+,/����B3"3cmhl:�ޅ������tx'�����f�A�������R9�N#s�c5��~���*X��s� m;��_m�9�AW����_5�l{�7�`b� d�
*�)�q;��_&{�$�����c˅�C��[�:}~3�w����-���G���j1�|�]�
� opD�P�"(�B� ���0dN�O�{����6��R�_�z�j=������|�����?g�뿿lrn�wT`�RRN�X�����+�<C��3��XA0��U���sW=/��G������� $L N�`�w��-߷��o��c��w�}^��ֲ����ѩ�S�`�?i�\�A�Tɫbo�2�� @�4 l��{��F+��&)�BV����@�\ņ��b�/������1��$�	 ×�#�o&=?;K�^�J�_����jj?s�6�ѥ��ܭ�n�^��76�rt� q�3%L�C����}|�$��局�.���Q���YA�ܖQ�(�����5�/#k��}�����(�x�̈́Y���;���S�߸�X:;��MN�ji~[�,2��i��آ�
8�1��<�Y�3�u���+w���x�O�P?��6~�I��7�����x4%�����jl��?�������^�)��6[�q�?�s�y�­��a{�\k�N	��湢U����|�+�&f�%j�c� %a[壛���[K�	+�e�U�ro'7/?>�F��N[3i3��v��tz�GN�*���к�tۭ���[��ϮItq`f��f�>�ߔKZ���n3��Ν˙�Ŗ�t.�ǅq�ѯ���v��6�r���ӟ�,��� �H�, �B  `����?b��?�`� ����X�Ϩ��y�d���>�d�0`M����;�#��|��}��$Ȉ�=^=���{Ҷ��=����g��m1��r!����b��D h]v�,�S�h-$]�O�~?��~�����h�揲��.����;f�ݧ�om�1��f��9������dk��f�(�f@�����u[ݿ��x+�������T��Lm��MN+��.����U(f �2Q���'��&Fd�ڞ���7�[��yg���='�i�o�!��=��ruSe��e$����kZ�n˛�Vy�M6���U�u�]ӯ��\�q�x�]��a���s�hd���N�Ĩ�R-˗f�IW.WNIE���
��,hl�d���9˻��y��^Kt���k}�)%��PnC�j��$�ᴼO{��6oũY f��G���G����cT�?c�}�P�x�Qt�Oߣ�&I?�ȕtBA=?s�w����_���y��ZR� ��<���q�}�۟���QDP�r��=I��7U,�J���i���z���m[���eΑ$�-��Χ�شa�g�d�r��;
��29�4 �Wh?;�O���0O��G_��J�H8�fb�������4�*dE1���H���]�kP�ddH�$ѥߝ�s�M���i[���1#'�o_�P��6h����E�S+����v�P�JU0a'z���F�ޫ�"Ĝ-"�20
J�h$}Z5��Q|������7���$ЅC4��'Q�<�S���DE�m�}�O�t��>D��l�8� &2;��$�H[���d�'��m��������ɦ��4�3e5��q�oQ�:�����׷��U����8::���}����"N!Q	��f.�7%Et!na����A���n77å:ϕ��a$4cP�k�P�j�OW4��B�u�.��̀����"p��̴���A�����'��%�q�0�ȅ���$|�b�r�-%�r+�^'A]v���Y�O��4KLd�.������,Z�4�ڒ� B�q�J�G���Qqb�H3��Z�z�����^#�|���ӌ`�s~mKh]I� ��׎�����*?T��R������7 >�ܐ+�m������g��Ta��Q�����;HCҀ��>{���Z˓�w���5lD"L��&̊+5�T�� X��Tj��(� ��f7����!�����?�
�A]�4@�2P���WCg�ax������!���b�g���0�;ݸ�j�;&l�k���Д�( h]m<��p��{Ng�~]!uQ�?�\�MW����r���R�W�AEq۔?r��~�(���I��=R ���۬����e���}h�� 2'T �1�P�%`��A����\`���<_9y�"n�*�	V��:;{��~<��!�b]����`�A�s8�F�/����?L�Yt�b��~� ��Eq//w���4U�uuv�g���]�����̋�,Ͳ��t�p���p���yp�H�3`F@��4���ݻ���9M��s��-ߟ��K���7�hS�Ey=~a0�%��Yf`���&'�;��f)�t�Ip �P�����5sN+� ���S%�ޔ��R2�yl���� n���?�A��ĭ�6榽U�Faԝ�@M0��r ��5�`%�0!0@I�2f+5z�qql�e~���C���6��N)�lDX�f��A��v#���FJ�'c �y�L�$'^��x�^2�R <W��-E�ep���_Y !��lbj"ߑ����n�Ap�B���3( �d�"c`	$MuU����+��讹�b��;7Rƚ1�``�/.��籫�`hfd]�̊@X	����:4�����5$��l���sIdv�?}�wX�$�'%��W�z�g�6Z�$�#�=^�X?��I�ӦI.���|0\�ܠ6�g��+e{����~��SF,�o���ȗ��Պ�X�D�n��������j�����c���t7���l�Vަ��� d� $<QG���t0 Ҁ�K��\�2�����~ 4D�%����r�a���K��=�=$�w9C]xo�?�����G��z���0MhH)�l���*�ڦ�I+�0/���;㏀]��n{��N������>c�-�� ��+i?��j�L1 RL}砷�>�f oI�en�՚�sj�oJ=�� ;���s��
^���7%�i��k\�| /C]�]	C�~�����@�X$��{����_09Ľ��?��cd� N�e��a��iQ`�N�OKg2�[�Ieq�;yv5�K�{�fx{�������h;����^����t?���On��[s�?���������~K�9bĔU����������-,�1	ю$�
�ܨؐP�l����� ��W��b�*�*<3�X�i4��-�D�R6{� ����i\RE~o����x��>?�-�V_��.j,S�g��6�ar��@��d���IB#!�KQd�]wsn�ƊwG9s*Cnu$��jŒN�.cR�.�$��[p�j6��ch�(�F��&��ة1�fR��F�	��������\�e𗧗�=;ӹ��I���^<V�5S �t�n:L��$$�D�i��5��cHh�J�AET���_""U�dU�˪�C�	RHH������REJj��4�[I���4!\�G#b���h�*�M�mB�V���?�I�*T��RB�*PQ��4�0j��6�n[x�i��������^f�j�+5���[�S�:\��1�wc�IN��k��7+���P[W�V�}�y5z"�GIwj.�wuݓ�w;��9�n(�nnqܻ�����勻�;�����Rc�ɮF��E��V��<׎������\����r�]ݮ���juR�軵ҙD(E�vSB2�Ddf���@��"��d_R�ޣ���kkx����  !i ��mC7�A����N����H��n�9F��H�mӣ̯O�Zg��#���g�s�$�Ԟ�Ο����R��#�4]�B��G����{[S�C�r�h-
�Kc�w��p��WGɼ�f�鍤���jS�U�i��t�J?�VbԨ���]�F�B�����F�l&B$$$hL���IhQ$�P���w������.;G�WU��%���N��Э$|c(���G�gM��I0�3��/�P�BV�ss�vGc$IA�[h3Pq��I��F�㴵c�i��.��sE��02ԅ��M��n�?���T�j���[5^�\5�n\��/]��5��r���US����8�v���9�9L4�T�Q)(�Q�%QEU�s�vH�s������5��s�s;���-a�ghI�9�m��!��}�/���xt�P�A�4�*�?���x��ʸ��o�w���U��|F��)F�T���CI&H��@�2�:m��m�Id���ą��r]��X��OV�(�"![q�z�E�4�h[u��m-��4���O�^&|D�.X�_堂�iڕq��Ȉ5T��*
�Zj�E�(2��*t��<�W��%m�rykH\]���x7`;,�[�͞��ǟdTp�viizUr�\�*,$<\ \��T�d��$!�S�6�r���Wa
v�BFRA�6�3 ε�.U* 7�\�UJ�T9e��/;H�+�&�:.CF�}�%��B�&���� Α޼8���\.
���:E�Z|�XU�w��L��J=!�����J��Ӫ�QTD��@�q�p��i�,uyG�vU���WH�4:HJ���4����۪/��2����pctu���f*�Z� ِR�˦q�
;�l�M��:b�Z7*�T��4�Z��V�$t����6�Ү�H�oU��"��t8u7{�Hb�,#d�*��jfofU^*5l�ʉJ�ee�>�q����\p�m}��2Ŭ�rY+&&둸#��Y"�0��J��%w*͡$�{u�U�k��s"��WJ�aLD�X��ʌf��B1��e��0�W�VY�YR`��X����w�k/i�e�]�]�TbgY5t�5*�p�V��B5`��(*� �N���<� ��G/
�Z)nTq ];�	����>��ׁRG~��t�R�����޵�E��u)�
utv�e+et��5-���P4��6�B� i��m�	n�zz��%ۮ�=�s���k��v���"�Gk5��Y|#��Za�������՘��(��8ަFAшac&8��b�Q5�%ѡqkz�V��RUJ����N���z��	.<.�N��C]�ұRcP���������#��m۸�v�OB��re�fL˷diD�^_ܯ��^o�̦����{w�,���GԦ+M�A��J��T�a�Y*�'��0x���6޿�%���qnu[�Vvq�.�ǚ�g>����β
Z�ߘŲUXW)"no��;f[�ʿ���~\��J7�'�S�M�hn{��Y���涹$����Dw>�l��o䳭*p;��u���(��Z�u0r󫿗?�t�'������6;.�wK��>{9�yO����_	�
Z���	e��QEWGvƿ�K���쓥�����\���2g!|j��J�U���Mr0,^ȌZr���D�б~�;c��s���T��s��d��`�7o����U�����wfG�e]���$�}�v�r��5�E�"T��Xer�W.d����x���\wck�w^|"��}��p�%�� P�m\�\~ߩ��@��ސ�E�C(F�۾( Sk�y�^ٷX-.(��I�f���v�Ѓt<��`����ヽ�f��tH�n��;���I	Cm���M�<U�%)^.j�U�^y��h�!�6=%�:N�T$��~μt}��м���{|�
\�x]��Ď4�J����I=��7�����=E`⋯�R���rw��y���Dss�4D�廗F����7���[���zwj-'7$\��{��߀����oW��}�{�q��љ����D��Ƞ~B�(�+�?�����	�z�Dt�%QS�??ԯr߅�$�]�C���[�u��Ýn\�6w\��`�w���͑��͋��{M_��{�r�x���Ik��xG����lw@?��9��Sq��
0�b�}��^��c��嵃8�
�'�Nv#�\۹˺��7���<��Qm*?��p�!��\~J��t�A!Einu��t��d/Ĵ}��������_��X�rY���~���V�x�`j��\h?rϖŚ��t��W����-Hp����Ԇ�R�~tp��F�c�J����]m������Q`g��Z�S_śN:R�n�v��g�M+������p1u��t[}N�X�f���ѝ�}�{ע�0�KnÎ�إL�eu�q�Q�*H�F)Ũ/�:���tg�H7���<�!$�6��}��"�2,�7���Bc*M��D��ImbF�R��	"T32 ��23`����W/�޻�;�����x9lK�߅@ͻ-��_��N�u�-�cN�ٛ5������P���@z�������p���+��	��;������6\��:,�	9jd.}�wzs7��N��Wj�̦&@2)�232G��g^QE����9�X�x&���Q�a�v��!���A`X�2��P�b_]���r�ޫ�"˙8x�D	��¶����lI�s��0{�#N�o-�_��ix6<y�,�����Z#5�Z�?7y�������#��[�e��9���}�N��e6ϑ�L�M~�����Ke0��
��]�)ɻ��9J;[1��+���oV���{��Ѭ�6���d}�R��k��)���f�?�R��e���}�:����c����/��(<|5ٿH�9tQ<ft�I'nuvg�u��g�w9C��t\���������[�i5���%�x�2�`�^ӹB\[M�=�3�7]nw6VI[L�Ѝ�!s��VY�'�2q�?f6+��o5���m�z��;��K]���|����U�crS-�����+1i��{���g�\1]���9�oN�35вB��6��s)G�9�=�7C6�v�̾�an�K��֎���z������fm9����D�ϓ�]�N��.��Do71��c,��{�m�[��[���g�P\��L�������Oг������pYׄ���Ohԧ�}�Lfn5_�������l�~��O������kd�����];�s����zŲmQћu�4���ɥ��������s���]�6��j�h�iI��ql�f�l����Y���cI�z����
i[�,������_va�=���>|��-�k�ػԷ7��i$�۴��5���]΁k&���֜nu�OS7 d	��� �M$+�ycT}��VUn�%� �-܋�@ch�{���qg:*J�D���7�������N`��_�t����<{v�o[Sk�w����Iq=��K�y�9v=�\Gk��ߝZ\5�z���C�~9g�\��ȭ���D�Җ<�5����=��O����/�������1��n����m�p�7��Z�M8�C{�<V��zs[�2q���� �||��a�7	)����k}t��q���9-��_^�4����N�蛅��;f���r1.=#d�GZ����'�l������'�ӝ��X���:�԰��djRb�IH���B�4��,�;Ot��Zc�-��}V"�)��..צ��tC����'[&��1AD�r����2�d����0�	��*�y.�{��j%��>f3���G&�$�y�k�}k/�$4�?Ѣ��/c��q
��ؙ��HB���s���j��ޟb)�?����M�M}�q��N�Ӡ�fPi�)�����6��P���H���R�N�E� �{��,��<wS��̑&D�	VI�$�A"_D�?��*���!x�}��X��r�=W��Af�P��Y���E����ؾ��?0t���\�B2��t�\��@���P
�&)&+�V�/R�����"�u!�^v�4�F�Blm�}����'��ǳ�_���|������{�qi�����?S.S�����s}v�5����#�����p.��O�u:�5y�y�iwG��'�u�
��|G2q���״�s�7��W����G��J�~&�huܛD�q�Os�ݺL�(��qׇ&��\4�k�U��A*�Rx�8�����8�%��`�Z�+���9x�/�l�'��=,���p�h�܋���:[�d~v�0e�g���Mq��w~dʻ���:�\�s�b��~��7H���z��_y�9�=��+q�xr�.4���@��$��Qp���}F��67��H���=��*��̆�Q�f�ز����9��`Ȧ-��%�莻����n���z�5ƨ,��D� X����m?���k����ĨjŨ��lfb�-�1_�B�W�*M!4����_ݩ�|�zړq�ƕ�$�U&䁙7��H#�.-	��D�=��9��Q..���G�/�
���ʟ2Ƽ,7B�y*��7��;>����v/����	���OKc$	������D!�o�v[����bB�������B�5��g�b��G�A*���������G�?7�M=E4�N_���f�����<���0 ��2KZ���Q��^_
����	n��H<��^��M��'�zy���b��(W������Zwx�h�B
�O��p[4��i4�Uۦ_k�r����&CcO���Kcs�@z���ڱ<��߷�� є�!L����4|��|]�"q��qhp���~e볚p�"��NN�����\K�Pe��i9���)�5D[� "�b���;Q�u��g�kKR��S�cK�'b�� �4�.�����C���� &_��"�����#�[_*d�/���n<��H�O�_����j��W��<x�έTa�@������[ոuq!��[�����o@_t}�\(���F'�|е��t�N5vƮ�1}��B��!.�e�
���F"���M�)~�g�JP� �Oa�&L� ���nB���D�-��) ������^�8��2t#E��:x�c�����ъg$@+/��^���c,B̝�>a^��AT�Vm���"�h�>��fV��	�0�ۢ�����jѐ�2KL<g��1%^Xy�2ݟ�ό������SÜe��ќ�@����ZP:�F	����]Wtú��/;��EDJ6��*�j�
���JU������lx���/u�'�qy2���A�c\�I�k���q6��ǁ���q?���}���@0�x޳_	�P �j*{�P5�xO�>�D�$�4�Bl3DӢ{��I![�]�K�Tj�BI%!m�����.@�~d�9"R���P'��nƚ�	!Xp��T�������l�Eq�������8X��t>ë�{�y��l�c\��ލ��!ű�`B�y��Z�x� Z-�:5��1n�)g�J�d�f�5D�}��=��׆"s������U���B�$�J����]%m�g�wI��p�⬟�>�I�zA��dKKn8�=�N�,?hL=Ya��>W��!}����Q� =}ϰ�q]��V;��k���f�5����~@���%����[egж-)���6�z,�I������[�������Ln�B���]7��~lr��bqDjL���(��?��Y�xpJ@������m��e��Lw��mZ%H[�n�o�aj���HF-�����,TDh�-��$)A�֯�S*mTb���0|������wx������;t����w<6�j�iS_�)\@<����@�ZT��ҭ*�bĒ�D��0V�/��n�G��qk�ZwYO�Ҹ�Ƣ
"���ҕ^�����ᵽ`.�R &���WM�]��.@�^9�GK�x��v`�Є�"�z���޻�S���Zޡ��-R�����#��Wh5�i�w�Q�ty 
���ࣼ���~O�zW$�,�"�!���5��o��"��K-p1�W��,Ml�r�^�j_-�˜\�ogU����zd�nC3��^:(�(�� �UPq]e.��;c�����i�;wPN»H7�"�^l�P�A��VQ�W .@1��v{_ϼ������>����W�KK�~C���eҊ��4��|�
���#��
��C��ܗBmZ �dn/[�nB9�j�B���:��F�~�@7� ��貂�="m|_h{�U�Ԓ:���E�ډ�!ţ�*Wg��*�+�\���꾅C�/~_L���N����=����n������� 5����/W�ɠBʾ-�<����;����k �XfF��$��3�w����hㄑF��(5������{��$�H���N�H�y������w�U%����yn��d��/*�)�(��O<M%�d�#&w\7v�1^w�t̙�$a�i5����{E���N\��R�5�K����		ی=ռ_˒��r&g���_Fh���6;���a�����P�6/$�y�i������.��ShY4a���+��}~~�M������7�B)�3�����X�j��={����J&h�N]��ei*����_S�i�\���m�_���F3H;��94j������$VA! ��*H��ɍ���խ֧�m�7�� Oؿ��"JP�,:��L�|�!�E�m�C Q8X�&NY����K���(H�H�F�[n�NL0T�S.$8�C���ruY{��bz�z{�D��^�) 5�Ly�a0��D��U�z.��E��osݽk�k�ԮE<r�_M����7���6�����c�6v�ұG�q�� ������"LA����ah��w'��F���%�g�@�4�j�g5��J q*� ��r������f\Y�,V�H(�ɤ� �@�Ƌ��^k��K���[�5�^��^w���Ӈ���O�^�&O/߼�����u�g:�/�.�9yޒ��ؑ�i\�y�/�G�^y��q<����@�T��E��\�y*{�$$f���CMCMv dt� pT:�����q�y�����HJ�T�Y	I�#�w�玶�HT���Ԫ�쫇w�_��ؑ�#S""�Z׽�շ���"i�vs8��*7x�})�d�0��S+ضȐ�%M6�A�<~C�Ҡ�z���eW�;G���a�b8�XL����/}������q�U�!���(��f�����C�󳎰m e�!5����P	(�"H�ܧj�ĝ�|j�:�L�Z��{Z�{��|?�=�\]}{O:v���l<�vư�6�RhʔUBU{x�u�v�6R�To�X�ɮ\�Vgn�\]�:չ��W�\�ͣr����1�*-E�nn�W@��FPDђI$$��1���h�� 4���zK�v�w��]�d�JwRx�#S�ރ=G��/�z?6���HFD4�<^q��
	��i`�ְ�'�C����~��ϳ��Q^�AT�T�l�Xl��r���ۃ�q�#�:1MR�t�L�Ԏ���ꪆ ��]ta�+>��u �R� @�@DLàW��@��;�y�yP��1��+�C�����0f@>G	�[Q�I.MJm9j��j��|	�	�Qj�N>��|>��ji�M\֯�w�sY�E��V4CJ:KUP�Gu��U����RɷV4���׾�<7_��VQ��[>vϛAw�z�(C�]�?"�4��#�.� 	§xq�܆L��d@�E?�/�]��ځ���Qa�Ԫ��0��m�_j��$$�^�2 8[��ӂd���ŰCd A�S|6�,�B�u��yCK�\���w;��Ԑ��j�4��t=?���T�8܊���L@z���I7���A�E��l��j"m�B���~��d-o�<$稨u���8��˂��+��=V��b�)�9W��s�y,F]�Ĺ/ʈ���/M���&�_S��w�l�mx�?!�
�"�i�i�bb"UUU$!ZN@�AjD-4B��X.̮U] @���ϔ�>�^�\٠�HYm5������]��z��vi(�#V�<C�J���۵k����*�wD�;�i�;��W
l".`�$�B"�*�q��t�wʵX]p����Й��ƭ R�p����H��w<�I`5�)[)R�5���.���[\�E��x�AA9��R�u�*�}�bAC��`�zz�e*>p�=E*�`�T<��*����T-<
�7ʣ[z����T����*��^�y�Eם �D�rw-1�`r�`(A�I�h��(�a�9��ܤ�7AR-�m^��n����������O����A�3l�l5�ȫ�*zǿ�b
��)�A�D'3�K�6��T�\{o���@�kPU#��_����1[^���K�222IJ��v+4�H=�:D���z�����w�/�O3���냘��ڎ\U@�񪒚Լ�V�{=;5�{'u ��J�rx;ӋC:� X�$Ae<J:Y{���J�;;���ŋ����������䆢D����;<�Ǌ��&n�h� ]���,D������n���j"jElm�@�	%���Mڇ������5�~&7�������o,��NʲeeM	0��UU��{��=Wd��;/^.� �q�z!�.E�v���U<<������GDI��y���
��Q�X�(rx��i$����3&+�e�m[j�jA������9�Q�X̥*oA��
�B�$��	T9.���<^�j�^�\*���W��-��$������@e{M]m��KH6��̺�ʯU۱ؤ�]��#�!���/0����	3����������	9ѫ�@Ҁ��4�WPȡ��|��PH)r�p&�so��_7s����m��m�#��	-n�e�����>�l�v
����=��o>�ODy�u�}^�U�*��s�(�4r��$dd$FDQ]2��!��peՠ�{Oվ'e|'�}_!�/�7j��l��iNã���7f��%��n��/�9'��9,]�D�Y%`]*�bĺ]�"m��}�(itAT�,�`b@�"q���m�G�i�>�LcH�B(�$)���@�?<��'\�J1D����w�����	S	�U9��<�U3��c�N��wz�9Q���*�04�Vb����g��.�0�Z��zF�Zr�)�lMlC�y�p s!�	r��7���BD4�k�9dъ\ZHh��.������ߐ�|�q̑���~_�V$��~�=��x>C�V/���@����v������;<N��?q�V%ђ���Z�yA�C�;��"��g��<��1Ĩcat~߀p���A��y3)����]u�*�C�58;���P�j�(,sx'����+��|F�1l�D��i������N��%� ���o���I>eW[�����& y
���O�
h����X�9߹���7�����C��2��5���2�����-oq�W�X\��?/ZZT�hS�E�4�TrC����>%19�)g�p��p�@do�B��g��������B��>6	P����>�5���Q���\yOcG�i�I'r0q������j$�~�9�_�p��~��E���'�T����	W�%����Q�Q�?�V½g��H�SO	�> �'����HOlSa3@1vTY�n:gR�+7�bg(����|�V����$e�)�M�[�F,[�~�������~��V�O���$�׍�/}Ą��hI-���f�o染	'�4�:q2A/�Q B��	�o]���"�����.����I!4o��=��*���>��*��I���ڭfpsq��'(`�la~J��A��.ccU����r�}zt;#��2�K�t\��y}X�7��:>���}���}�9������ڇH���۴��6�#>h| ���k��w�~����yW����_o��;r�Ƅz���f�BG�x|6X¼�A}1�`H��۪��!^�k׳H���X�M������^�\�� �G+��Ӫ������́��wtЩ��{��h�'�!=t��0T!���Ţ��ȸUV�r�Ț��+�!������Yu%\�B���Ɨ��l ���2�o��C,��%��b�Ļ�^?�h]����{���WA�quD��>���#	J���@��}�����]�yk��3]��W朩9"�2aM��h��}0��`ИD�\֪�tK���FB�t9��	BA�qKB�V򭠟��G49����n�`"a�3��{l�A�1Up����=:�K۪zb��jM;=_�� 8#@W���H���w�[^���=�������8�[�{�R�}P�CU4����!�ﰪvU��ep!�<�Q�
�ϸ��S�^��W!�/iA��eTD<�����W��9�>�����?u"hC.������m]��c���:�h}^w��ݠ�)'���I/��NgΔ�������݌��T�*6�Qij�/��M�?���\>��}�3�kQ�qX�O��[���=� Q��3����>������}��j��B��X��*��lr��bnh���9��a�G�~�-���.���k�o��A�3>"���BI�!*�Lqj2�ͨ���m�ڋW���{4�BBBU�l*�4���{s}qO���gL�9	���^�gG���Wa�)�-E0�Yj�IhZ�`�[�L�gR5`�PX���v���/�'���k�B`;x]H��z�<*�C�!G������4�*C�JԑD��y�+H�z��kt��B��!�~��Ϳ�z���"U�)��-�ϗG�T�� w�tf0�}��7���+u�ic�k����bb�TVƏ%��1|�+�UVH�]t˷����S�E0�D��8U1	~ԷymgZ$�#|8H���?5u��I��ǒ�Ѝ�&A�4��N���z�uY^N�f�	�����e��\c�q����t�p!�>�Z;�W�bq�,����4���_6Ťr�g�9�<�B0nω�&Z$a$$/���Լ��)�p����?z�i*6�C��s���US�&���r3�hq2�,�j5`��mRY�p���aRp��?	��l��T���f��Y�q A������6e�T�#���^f51<��J�����mD������@��Pt��@��M�ibW��i�T��υ���������2���!hSƗ�>�K����!PAg�����SK׵��/�?\ߘ���BjV�����H�	�8iT���b���`�7�gɿ��>�}X�fI����>��!�����%�+�'���o<�h��:��3�����t��|uw������������G7p�^�I,�HX��l�B]j�U�=�w��w��������=�?bC4p��~�^����B�/�H��;�$�j��-D�\�1s7��y��vLX��]w1�K~�7�Ld9.�%��*��5��ʷT
�W�q�����|r�"�R��U��Tq������,��"u���'��I1s�j�p�X�/�y_����˧p%k�{���}�yC'�V�k��#y���-y?�b�(�<�VL^G"⹾d3��q���v+������ʋ����G}���vR~�߫�4����=WA$��`8k��D�����a��3���]9b��rEš���g_}#j�W�ξ��@�id�T�(̳4K�͈ب$���������������*@j%��e~W���!$q��p i���2���M,�2!�v
�c�ҷA��	�5���>I��¿:���\��YD�������mD�����.{UJ��ڣ��H�Z�_�@�Ef���� Q��F%F��X�>�KEj�@(����a!w��/�r�R ͒I4�O�W������>��t�9\1�̦��̆���`�zn��bB�������O�CJc��iR�����|��x��i��/�����~��ba7�#mG��>�s��Bª�М����a̚���D#��L�g��OAvD'�wI���?G��o�Ve~��Jo�v^��p�Q�2��[����^�äzO��c���r��{�~�Q�UC��
��g��G�$i �r09U��K�/�,��w�Z�'�Ly"�N$����¤p��h��m���C!�,�c"�0v�ƍ���^繢�G��M!��z2�tN�Z��$1��>��p�_ŝkVE���P.�4��m	�����K�J�3,.��So�o�v)T��9� k$#dlH�$t�$pcN�Q1}��Q��-"c 7��ld�qr(H��� �\m(�'�j��x��2	 	 Ȅ�dٴ_,ƴ�i��0���߈�`���������M�#�ο���=v�;v����<�p��Iqx�`ैe(�]>g	��?��5�b�@�a�f�Ƌ'j�8x� �`�H>�6Y%��_s��~cȝ��s�3����7�j��u�*�e�3EVeJڅ�f����5Kj�Dlmj5j6ح����	mf�M��mFd���+d6	���6���lem�[J���Yj5)fU���hM���[If#j�j����6��J���������Kdح�`�j�QZ����llj�Uh�V��Z�j�h�b5QV*�Fd�R��6&�H�j�I[F�6Ţ6�h@I��j�[����ϟ��H��8�M�:���ұ0����^�_PF�Dd���@�BEޯO_~�����u꽿�oa.�/�����p�ӫ/����o�zb�HS&J�W��?Ns�<�����+s��6�>��!�M_�s�	>r�$�5}�b���1?�-9\P���0�����c�w�9��|���=�/�t[��5F�j*>7�������v1{<��TՀQ�a�����>JŖ�߇�4�0.�P��R
!#RR5�t�w6ۛ\
��Y`ٛ6�����-\���+��:�v���sss��[]-�-�ssd�������ܭ�������9��K�Vj��Q�Cjm-�ڒ��Q��M�ء��`�Ҩ[QKhR����ElH�ڤUl�E9�̥G4JfI6��H捤F�֭���r�#QW7-TU�k�-sW4Qk;����ʼм�d��i��*��4i(�lX�[$kF�-�H�5�ؒ�+������]N�r���ƴlcEnk��6��3XأQcX���V����X�&ѶJ�b6�Lbō�b�IJ%��wk�-��h�Z�`����h�j�w65wv�TZ6��něA���<��|��~��T4��y9~y-n���\�9�<��:����2^��o����j�j������o�:�ߏ��v�����?�f��i��­�9��k2��Qm �3�̓\CJw]�;��,W99q�p��#ݮW3�cmnI4�j��k��bl6	J*Qm;q�F��clI�I��3[\��̶���J�㜶��]�ӥ�"Z�+��k�l�cm�6�湕����5�Z������sDo;�Z��\���b��f���ک6��PB[6���jlm[
)[F�J�emJ�m$�QV�Sb��J���m����jUM�*�DlB6�d ؕ6�F�"�Jl�$&Ж�)m(+h�6I-����m*��U���Ȫ����*l�[ؔ�E��L�l��[+���Tڌ����ѦM��b�7�4d�̚mD�wt��wvX��w(��dP'5̔I��s$�) �4�j�\�;��m���+��ɉ&�Y�W����U��\a�%������vr�Q LJ�@+�gѢ�R:J.�������F�I��o����~�=M�c��j�z�����y}oEU��Nv�-5���?�����zuq;���h�Zm]L]F��G����7��G.��a7Q_��'	GU����Y`���k�����q�`�~��^_���_�ŷ�����Zi�1�A��Q�
h���j12���iqwv鄈�9ݮ`���̬�Ri�E�r�9�!#�sH�$C0;�n��:pNnQ�ΒI6��&����4�(��(�FI�R%"�dDI�0h"$c"S��$b	�7]Ӻ���()1��]� ۻ�ۮ�i�(�Ә�]:9�5٤2L�tƒ1&B@��%"��:�ѢRwvE���n���t�B�r�	�3�wI���f	��)���Ąx�I�I��$̑���S6�苻pa&A�FhHH�"L��$�f0(�%�s,�a")Wqt�L������#��;��&F�aR]�"�F"��ۻ���;�Wu�)�S�����';���w\g���1L�L���@�7w&��hJ�H���J�G]v����"ʋ��w�4JnvEk�Q���wWyܐ�Q��)0�Ew]�6P��.��2��Δf�	rD�D��$�u�2A�]�5�wq�H�H�뮹)��bR&�h����$fR�)i�2h�.r(]]⻝��t�tݺ��/���� ��#2 _�M��9��c�w/�7�Wg#e��}��;�_�<��O��h��L'�a� ��>������k���s��,̧�c^�)A��x�߫�+�r��l�kd��%�wG����1��܂�X��6���v���pN��9����9��+8��k�����}���K�]���m�������rO���i|6�}�J�^v*�e]��v��'4OKJ8��a ��	�aj	�&8b��H�QA�-$Do��L �"]*!�+|j+h8���4Q�b�+h�6� ��ⵅ-�K�Kaf�FAJ�4P5���+�P�O�DA�*�E1�W^�#�N�]hu��ݤx�M�Y-*����U9�"�Ȳ.ѵU��i':�]F��s
WZH>3*�2*_�D��Px�H�d�ڢ�WY	]`�s6D�H��u���EU�IS��*�"'1B���sR!�R�JU̥#h�����T;n`[*�(��T���J�`B�Ul � �$�P�ب]iGl��O��:<U
�%ҫU��m��N�r��\ԉ�]�xwp��,�=;j�d��l�ɐsWmO����ǒ���ɑ;i;���ߤ���Ư*���^�ӬwcŢ��ߊl'm%Uh�����b��(�sςQ��q�q����E���qކ��|��T�	�T���UA�0,����æO�������(+$�k2�o6@��������������������������������������� ��{�t ��T�       4h ��  }    ��6C��->�QR�$��@�   �%{� H� �|n.�@|��p�(�`0O<�qR  ;[�מ<����x1�{�-0�� ��{�<�wA�ѷj�t(��;�g�{Ϯ����v��{�      =����=�޹��o{�l|�D     ��d�@�|  ���+QE� 9ݷ4  �v   �uu�'bJ��P ���
$ �- >h��a�5�v���ѥ�����j��B���>��@G��� �\��7O�����e^�0 @�<{@  p�      ��x
R� ����  M    �d  �	�F	�����Si���dhe6�hi�c�0��2�45O�z&1Pj`&H@@�&L�h��S�i�4 � z�OQ�CL�F�  @   �!��d�d�@4S�"HDHyL���!#C@ z@mF� i��@ �h4     P    � �h�IꔥG��444��m&��#���A�@ hd���� ��� @��d    4z� ���jiO���y1'���zC�zz�����S=��=M<�&��MS�mF��4�M���a4z� @4Pi� �H�d4i�@�6��OѦS�4��i���F&�4��#@ɐi=1�)��1&��&h�MO	0�M��54�!'�&�w����b��P��p��g�{n��IL�|�#��f������廻�.��n��fm.Zm��ni%�B#$�2�w5�\��&ro5�UKd�Gxn��/c����s��e.���<���g�������̃R�1"Y7I��J%���7,��w:w�N=��4��8���/7%7�t�!P���ݫ�r*��ͼۯ����fC�-\�c�K�n�y	˰XTO.�rNC\(�"yCg8M��4�&���ޜ�kkݼ����N���/{��_�;\yn�M�*|VOfQ��sJ2<�U��S�7��z�����$��p���4Or����{7�\����t'�1��yV�!'$X��
�6�a���<�lU/l�^��ض��i�*���=��
�������>D��>�Ϧ��fšhb���B@B_u���P�~��D�qb���|��~E+� l{$I�HB��Ȭ0g�\�t7[��r��`�Ni��Cu���%S		MHL�1�2���}�D�P&nl$֡��Y�L��n����2K3(��53������%�Wt
fd�a: >\ɕq_�ߜ�3r���`.��*)R�E�:���J����6�I�׎߲��v.c}�{׸^׃�5�^��P	��e�M��;0�@�xChdA��Fp��O���TW�h��������x����M��q��?��.w��� �ID�@"�f��r������*�
"�2\�R�l��Z��	�4
�.����U��B�pД�c>���p�-kX ,8��XV�F��q������}�UH�h�́j��w2\o����Od2��e��5�nS#)�1Ҳ���B���R�s���L�Ң�������-�֋r@�VB����E��۞����v@cqk���rknQ���WGA�xu�&ձr}Mk�i�"�G�X�dC0�M|�4�u7��F����&�|�s�ӫ�fZ%��y�R+����Ax5yd�4 k/��o�"� 3�-t :�����g5��\���IP-�,���#e䙖q*��L����d��b
TA��Չ���H�tty��VD# ��0�ƃ�)$%�0�"+Q\�Dc ��Q2N�
ąa��K	(��@`@�#!��8�'�lH ��7�p࣓R����G$�ml�����,�v��S95�W��,�4�֭h�r�ӑ��',8��Ր(gAF����3#[l��!2��V6�;ܒ2d�<�K²������gsmtI,�b�p�Ͱ�\Au?�d�� !ae�*��H龃K�N6qǈ�+-ۘ�n$P� {3�/	q:I>�)�%ĦH1���²F�Ƭ����b�es*(��h8��St�<�)�ա�L���d@>PgLG��^�@<�^za.�| ���'���"�����R ��^�̬E1���|��)"�J$�#*EL��֤��.޹M~���5�]�>��Q��_��݂T{f������]��ar�\f��W�f.LDE��A��y�{�l:�oæ��;z9~S�sϠ3˷��*�[B{��[���b�������'��;u]B�.Ene��۸-z[�1)6D	#�`�6(`����Ux҅F�G�p
9�b@�����@��}���#t�%�M>�
����D	,��9.0fTWa�zK�;GE3�z �H8�s6�bۇ�9��R�}�=���َ�4d0��v��ݩۻ�y��=�M`G����+mN�Å�^|%�)d4��x�=J������a�W+?x�y�(�����}����Ќ/!��
ݜ)s&)�=�OQۺ>a��5� ;˻�@��x�z���{X���
@T� �����6[ �c��6R�)�:��]��O.Bݿ�����'��V�o�͓��C{׷�� �nOa�p*��H��]ir��pl d�S	�l���O���UH-�Y@��n�Q��p	n<�ɡ�Hԧ�%d���b���������,��5�w[R�n�I�n�:�_O����;��ȻƧ��#�8�GL�>�S�dL0�z{r>[�l�At�[1��g�zן�M��;^���~d9=W�j��~:�`O-�}k�>>��Ѿ�5�����.���}�k��>�﹉ϗI�|�m�o��y��n>֔�۹��k�0�L��4�2�%�3�+�|�5ѳ=*�G�6�g���mt��mi�5��cF�H
ȱ�ہB�b�`�/�E"sָWO���Ғ%8���q��}w������9Ws�2�=o.��zx�h�u��<>�g)�C��^2y��p㋪�9�$c����Z_��ҝ���ہ�|	wU�,�Tg�mT>�\�]�3��^w��3K��Wg@���S�%x'L�9�%e��WB�fκ�d�e˗�~Y"��	�tþ��o�=ͺm ����%$��~�Gǔ*��8pP^��u�{�4۵�u�Ei�u���t�i됊ӟ.����s ��c�]����4�S��ɪ#r��܉�j����oL^����z�ɦ��_r�y.?K�E��E$���=��o�n%t�B{\�I/���7�m�P�u━	�������:���חT������r��N��������˶`��;��zf��p���]/Sc/W�O>�ĺ�g�
�o$��e�yᷔ�2wl���Q�:wji
h4��5:�"]�۾5V���+�z�-}<���w=�m�������nU�<g�6YsM���i�d��ǹY�^���o�-�%�j�F���`���)��da��}6'���M�2zd[K�n��g^R�e�������W��w�i���2^��d�r�m��\���_�.������,	���<���,J!l}ӻ��|c��鈉M�~�>�x���
�5:��ݼtG�0�gÖ�����lVO��t���F��ee���ɍ_~����BvU�7�>��=��_^���o�ڍ߇w����3�ᆛ�l�k�&��7�o���I�c\-.�_1:��ӏ�oZ��-�htt�	�#�\������y�챙�l'�_<��um}x�uN�Тy']z���g�y�!(S��s*��\J|o���ʌ��k �6�>kuR7���&��#^T�̱�	�~�\�=2~���G�C`s�8]�/�7e�]
.S;/m_B�˞m2ұ�|����8<&��>x9%�舴��ª戉�pՐ�](cl�4:=��JZ�A����IO�e�Z8���{��Z�5A,r�Y��}t����i�Z��;����Rx�n��&$]3���>�r�}^���ķ#e���s�����g�ۑi��}�\�[��D�Ynגޏ׳�8�L�d������<���s��φ�?;��~�}��E��z�=Bj1�9���LL|<A']_1�L�+��IWi�7f�K���Я�[h��kQ�������ׯ����.z�˖���/�������:��m4Ѡ������}���k��.�>���ȹqR�è�� �ۍ������k-��kE�=�n�6��	iL	�܍NQ���$2�9)OEU4,04W�g*��!�*�!���$eh4�]�:ʰC�1J��8w<D6ML��t�?�|�pV �g�d�@>x��~\�?N|@�|�OlƂ	��A[<��S����nn����5�0�U�5�¨W0Lӆ&�Ec؝�J��ҜS(G5��7c8$!�g����ꉬ2��з���y���H^Q�D�o|���+{o�^��V�w�k�!��7� pTn��2�Bȵ3f3d����s�0'��$��c6"U8\R;�1�
@����P�4�둏Onߪ�"��Ϛ������k�AtHX�4�h�+a�0�4����Ȣ����oX�،:��Ζ���8�0V����m�
2���H�hh���G)|1�%5*�f�G�����uF?b`�AF	�y��K#�>�
ml�uܢ�Pc2�F(Q�X�l��� ����Y^c�8]�2f	��x k_�>E�R�(��{+���%Pn4ՁF�c�Ƙ���<z@���Yu㫏ӠL���NCz��Ntr�\���� 0;�$]p���	�wd\����H%lh�QA�k��a��/�A��Օ@�P�5��5f����!«1�ō���YS&�	��lK�K�R�^Kq3&������"���ۣn�g���3M��$p�3��/>�2{�F�Z���8�B6����LH�#�ma�� ~��/ÿN��{s�.��vӭ�r���m�j�|���{7 E��4ˊ�Ԭ���La���M�Jl�^ܼ�=��2���Zs��Z���˩�U�ɟ!����O�#��HԏG�"l#գ��lŠ*T$:�1A{@�e�OF'�6X+l�(c$q�����Xa���5��F8�p�8+_�:]�^��jI��/K�9��FN�r�{G�B�"$�CVZ�h���3O��&�s��6j� ����}��Z���|Wx�Mx�6.#����]<{���c=�ܹx�e�Omdxu)A�ۿ�|;���^�S�h97Tv �I��RĈ�|��<9-p)�b�h��CK�. ��Aq0��~�/��[t�����{��:����?V��A�[�c�`����J�af�,�_U� @�+�F�|P\!	叅Q�v]���3ڱ�Hm)
_�SS�����<�]�ر�wca��;?��!�w=O(y��;�	y�fpҫ���uS�;T�t�̪?aTY�+:T�̝�M��/�!=��/�,�C-˂��P�C� "H��B|e���@��N{p��o����X�'������߿��Pڍk;�Ŕi��TA���ӝ�Ȟ�mZTz�w�PE<��Q�?)o�0��d��r��SK{c��m�'z��i	5�=9V�V�{�:A�@��U����DnIqL���I��ǻޟ`Iȋ��,Ă9{&pO܄|�8mq�/ /��M8S������aQ0�Y�u�BVĦPQqM��f�8�����Z�L6�X�7:���c�llMfjDTG�rh!���7��ٴ�Ò������MJl�77^�,L�]llv&�p��0�UQ�&��CEل.L XS"9��5�t�i�0�g	X���q��
L�\!I0��J�ԙ����ɘ�b��9�&	�2H�`��a�7��)��X�g5��a��S�-mr��ɘ��g0!A;9��\�;w������u�b�"��U];��\�:L��9�I&�k�ٜ�q)91�yw!�n��nf�	2�����rv^rql%6Ŷ�˼;������y��w�y�ݚަ�ޗ��$^��[ӗyq�n��;� ���� MC�hW�<�"��XC���7��g,�N�vsy���+�G��-�y˩	l�]4�[ˌ�,��&��<H�K9�Qh�9���w��u8q��Y�9�m�-�k�9g�6�S��^�%�D���^�6[N�:�o;���צ��w��;�^�G������diyyku�����sY���쫽[�[�Լ�ڇ;�y�]�὜���R�{�z�zi��'E'/Y�7g{6w�'^;�ɢ��5X�Kɧ���f�z����/+��n�UlW�=8���,�x�R�-������xI�[�vr^E$��N��D�^�t��yƥ���lH��vF�X�w���wk�qJ�Tׅ;���ٲ��xăӗ�Խ���9��p��&�y�&u�:������ꝇ!�d;�����r�:0y����ݛ`.�n�Y�N��u�8�����\w���x��8L�P�����K݆�.���E+�yBH�u݄we��D�'<s�d$�rE�ݧ8��lyhp�s�ӛ�gf�͔J���#��{���H�{�Ey|�<��;�7���:C���;��)ÝǷ9����`�h�{��o7�eίv�,9��\k:�9���Ν�9R���쳓�t�aNL�/)8�Ԑ��/joQ��e]��9oN��&����פ�$z͐�s�{7s`�m���u����*�N�(j��� *
?�k�S���G�8�D���n��-�jME��*2V���#h�T[�E��Eh��F�5>����=]mVdl���l���ϫ�����Q���*5[�&Jɤ#)s(͇Ezn^�͂ �����v�q����}_��?+ۺx�*m�L�4ЍZ�1���1P��SZJf�2�%��!OWD�/���������<��[ �S(�__�h����+����a�4Yja	A�B1��i�.����t���03E��Q�Wߍ��,��Fi24Y��v<�1H,�^�����Ն5i��$H�{����c�r0hrv���Y6�ܰ�EdK�
_q�`�d���+�� ��VD�ݯ�����5����9�4��ѥ�8�F�4&�M	��U�c�
t�X�Tǈ
|.�����΂l)��1�g�} �o^ڨ�G?�����u���?5Qyx����3�������'�껾��Rwe��%��(k�y�u}��3��9ˇv�ke��]+ ���������^�w�߉a�|w�6`y�z�vq�1^�_WO�٪l��rgv���bL�>l^]��w�R&�iQ5�O�P��YEa�m�kNf��A������h��+[;csss��isjxnen6�l�������a�ҟ��b�F81it����r��l<]�ϳ���{�G��O���\̽S���ػk5�lU�j��f����y�܉����x�g�`���P �f��y���[q�7+��x��  �@���u��[ʏ���9����pۉOZ�m
�<I~Gw��)�՟�پoX�]�u/���m�{��<���s�>�m�Q����3v���]���66�Y�+����r�Y��&�,9����]{��cC���x��7��VڮΥ�5ܝ��4���uqj�i���\U�Z�Y�Q*̰js��ni���g���$�޿h������Y�f�u�������<�_`�N>m��*��j�:ɺ�������G���kr7C�&�o��7��#���u��Α���3/I��Z�<g��7�a���8�n�28�?5l+�+����o6%p��`!  �0��z�67��E辝�Ǆ�z�Y�3�!Qq�!%o�4�~��UX@8Ҏ5T�0��fpZj��=�m�(Uh��wmF�'6h}���Hfi�D�z}��g���j�;/���9�m���`¦��U�O�{�m�`v֯�����du�S����@ � *��
�NH�s��"P���" w��E�G�� �B��t7�'ǐ�  21`�&�QX��js��1�7�p#�hf@��*��hr/BU�����Bxȩ�0�P6� .;Q�QQ��h��S'��t��;O׀  ���H!("��k@��A%6aB<&E��k��4��E] !
����r�w[
.���d� 2�n�A�r�?9_�������XX7?����d��鹿�û�}ȑ����tNXj�N�!'�<��ƌT��.o�Ȅ���vF�s��$F�YEB��# bk�]J�R|#��X͟>�*` �|�t%��J ?�er��̼�  �E��T�)�z�|F�ٻ]IG)/y'~ � 	F�N��0�"�K"�B	t� �-������xݱaQ	�<�T.�;��?/�>��Y����X{, ��w�]{��!��ܯ/g�S�N�zhJO�>Vg]��m��Q_��G�:w����w嘏��6�<�'�6%@,1���3mHU��,����V9�W�"�Z1R�} �����~Zg��|N��k����wŦ�� E_cf�_��b�`��Jc�}I� Z� A�N������c Ye9�%�x����_��Cl������_.<]�u"u�n �|�}��<}t�-VJ%��`H�!�B �1 Y�{Ơt�
��l���-��eY0�.�i�y�(��ƛ�mlW��A,C��@u�"%b��RE:I"��1s������R�QYf���{��2����x����1���ֵ�?�����n���&Zz<~��i���;'�w���> }6��VX>i�~�{���T}K�)�����F$y"O�< ,�@ #�Q�M�`�qd�P�vʪ�@Y�n�2h���X�+�*�j�c'8�p�5b�[��(� �^�Ri���5�*�>�_�:��6S�!ڀ�J�(�>)�JÌ`_в��Sz���ƪ�8�qZS=}u�' B+��Q��`1�
Ǡ􄲞{�^!�K$�ܸk�C|�4P�qe�1���H���V���4@ L�p+FU���|3����ti�jd �d����A 62DyLed��a|�lĚ GF��UV'K�C2�Y�G*������B�m�]�uCN�И"�C۟1�"s'�4,n��q�<|��4!Y @u"
%[�! �1��+�����D��/ � ����v��e��c�c�3F���fOj` ~%eaOKD�H"/���[��F��Y��iƙ��I���-(�G�B�u�5��	GV#���Q��W����?��>� �ak}\��N
z��s���������}
<d8}�e�O��<֜�O/�Ľ���B���0AI#� �r�I�v�n�μ�y�P���Byf�q���J���,V2��b�"܈�Zǂ.N�c=\�FX@  >crM��ud=�5���\����̓����AA���L6��̭LV3��c#�Ά=N�s�]~X�o�_G3_�ׯo�ox {�����сt�*{�����}���qӔnH3cT�
mEo �)��T>������S#�h&�5r�L�8� a�l�jE�e����u����SU�x�:���^�V��$��@�@߯0��D�Ɛ��N��&D1��v�4��ʆP�1�v	8�0իATAL  IKM)B(:��0T�p)�4sw[m �0C0�v�xe� f�#t�@i|����` D�8��M�7�o�-`?"V 3�_��}5q��t-�8_��Ι
%(�͆�|��%�Aڬ9�Ż$B���eo�^�֓|������C&z(ʁc�0�)R�v�6u�
=L@���h�w/w������<;�a���y���~�Tc�0d1�GEr�<V����_/��ehȊ��#"��F�:��r&d�KA�a�{���"���/�V%>
��@��詝2|ʤ��"*�  +�~y���pB
u@�<��x��&|�s���XR-��(�5>� ���.�Fp��Ŗ1 �M�ϘjDuZ� �OCU2�[�+�
�Ą��e�P���b#γ��C]�A�iZ2�D�( )��t���w��N�(��b ��l�+=WG�u\���:̊�+S�,�!�G�f\3�R�����R�9��6�MC�:�e��!��c�q$Ѿ��s!H�i!�5Wt�9ⴌREYA&y�r�� ?Vvq@�t����i�����t�5Zv���D��O�@fd��d��#��p���@ �����!T�bZr�MU�������ttѕ~���Ea�D��D�C]�2Dk�D�F�~(�e�w�~H^fcq�m�ً�fLb��A \9�Z�h"�Y��#�U�f��٧9��%T
��I��H~��X?{{,����XH�3�0�9EXq���2R�S(�k�~�.���*Q��
h��Z@RiOp *s�bY	�@MbP�s/A��&�'��[�R�H$���*�j�92��a�x���C�!&�gXA�����ͼ�;ϗ����ަo���1}���|�ӛ�yH�ʬL�9���)�T04u[chA� 	 ��y���G��ju�	b=$]�:��2i���+5F��U�� �:���,pP�Y�����@  ���*Z�&x��J3F���##AY��RO �`\9|�qIr�Ta �3cUya?�Fi9����ˋ�-�&��EЃ������HhU�Tь��܀ 7j9.&���RǐRO���3rxYP�U^.z���]��|�Sa�h��U�[��6��v����,�1j�r��i0�C]�k벺�J+*7�T�����r��,S�IZ	��3"՘�wm��eB�!��Bj;R�`���V��	�d�H��킩&r�.߼�a3��Ʃ�ݽ7&��D"(Ak6������gU�Aw��c�mK�*�Pu���n�0�jj��DB��9̨�jQ2�4ȳ��,�]*FU�Lb��͢�t
��@)� z:�EY���oD�1��ϧfV�篂+���C��,��� �hdd�3�@!]	�-�I
V�cP�@ ~th7	@��d��@�0i ��@��sw\p!�&z`�2��*d�7~L*-p��pr�B����L�<&��e�JB11�* B->B�'��;e�,�ԉvd�0@����NDl-�p�("d�a�����u�B(��	%g+GFŰ{�( 1I>߇�v�=��q�3�f�a��������ʞ�Z�k�h��lK2  ��@�ځ���Y�k�4��(� f!�֏O��١"��b���X��F@B�t <@( @�\�{�33��5	aEi���P�>���
6�R`�摈V�6_a�,,$C  �gf����6������I:(�Ip�-H^-\:��h��@K5�E��E4x�����l��l��c��lX2[/IA�q�:�o"��F��8Y��Z�-�$�Y�o�}���6�g1<*N�q�B :8�<bx�ʈ�$׋���䬬
;&2��,�����;���P�ލ��k����+�[O��؍\�c��w�F�ֿ�H^%�E��� [�,>�Z϶��l�ܾ?<���և~�D(IЬ�:�ܢ�ʤ40�@�X�5(�akZ�W��~~4��xr������K_�^��i�.������x�w�鄊jI�W���["|�����r˲��07���V�l������or�����æp��whᱴ׼����tr*��E�.����V3�F�d�[FB/	"v�&�l����9I]�MMW�[o�������S:��H�N1�9��7M�֫�s�Q�Ðg[-��wG���ɥeͲ�p��hSe�h�\�C�
��@���b������V�����y$H<Y-�`7��kz�Y\�.��!���#�o��y�5�eJ�o7[�ǯa&��+�rA9�]� �B"���{z�;�3wzvt�#�w�@��YR��6P�׀�מU$G����ux�����ɹ���{�-h�����u�8�dm�Yl�ev9�'$��q{��y��weZ��[J"ܝn���):��6�Nmm�C��b"�G9,��3f����p��N1��ӗF�Hr�Z��9�^���Yh� �����ș&M�KSK&�U��j�MH�����e�ja�L�w_.A;��a9�S`���v�ް�6s�C�jIĤfWX�����;{؇ �2J�Y5���u%ć�X��+"��R�*���U�3��KY��a(ȇ��!�3nFY�8�\Jҕ0���/6�)"9��d�^i��j��`��V��l*�ؚ��;i),D�W)8�M�RE�4�3�����T��&9�ZF$��1�,yFrJ"��ۺXM�3�.��Br�&�*Ykgw�N$WL*kfr�*���8�e�Y.�wdnL+i3m(�[URvթ$W�7��I�Ja#�YKG�v�J�T]�NB�5p�Y	�+�YI��4�,k�8˰��\�,���u��d��I�X�8�����^��ֳ�%�mdE24�jW�j�Q+�F�-M؍iI)��������b!� D�D���R�����O�i��n7jN48�ƋcqĎU#��<�6�^߱����l���Q�Z��5�k�,F�kb(����XՈ�6��sTb��V�`X +������(�j��j�.��� Z���ZT�+yC�]����'8����<��s5J���Ju;m'g��R#뻶�$�s��LS�7o�=��c�����lTbƾ� C$"�5i�b�i�z����ϛ�?]���v�<�Y����螾M�a�X(�F��P��f�iJLh���FJ�$��@Q��h)�dHERBCL��l�$T��2L̊�JMȕE��X�Q��cQI�e��EDl�h���@
@b$�EBY��lb��$�H)'G��y����:G����䭞8!��3����mi�]���j�H�(�e)Dm�,T�4&��d�5kPQ�#b�bA�d��Q*���F0���c`ƣld��l��[W���.��.� B&+�y��?7���?���"S����Yp��/�P���V瓪�
�k(�m@�Ac���g�s���L5g�96�/ۂ��~>�(�I���rwO0�e��P�����:(U�,��qZ+�+QCݖ���4�S@eVL���Z��'�J|�>~,�e3eŖ�#�)SWY���!�ݷ�֖t���է�v��5V�[n�፣p�-Jyx  ��������a]iouE�P!�j�%��]�R�ą���5T��ŏ�nP�a�T)�"��ܫ/�����u��a��y����?9�u��:�6��}/���;�N���~	�%����'~w�-yZ�RK�X�12qI���\�9}�Xȗ����uu�&��dH�"���̮�`K��\���T��b�0΁��[�}����Z��������_�p���n�o~]�K�m{׶��;2=rC9孤�нE�l���8�E��= ��/�
w��6�����L��w���
N�H�-`�
��"�e��q$�?ϯm���({Z����:�ySMk�� �QdK��9��o�VM�|	����/&TtºjJ�N��u�~������<8s����h[+*��a樐��Q��f��D�ݻ���F�����i��CF&2Xؠ�`ƴ`�,Ѷ�4�)"*h��cF#d�lZ"�
TȎ,"2 �-@VdP-�v��&^�O�=ϋ�?)|"�}�*�����M����8'+����e�Wg��Wv�t�(N��]�J��^l�͐6��a=�6�s����:����p�)K\�R��QM�#s��Z��)l��K������=����J��6�c�Um(z�a�q�L����XQÌ�L�3"��`zk�ja�b�����/�*�����GO�H��{�ڼ+
0�>_3����`O�]��8���{� �9����=�������~|��`�0s�=�e��tvpU�  �
~5��������i#�B ��~5��B���J*	 �I�N������n`%=���@��7�)}���F�h#J�9��x	ާ�KJR���)< �B xo�����ԏ��n)K@՟�j=�O����z>x��U�(����2- ���O��t�I���+?�Ϻ�����{�У�撪���i�l���L}914 ��H� !�0-���.P�Q��")�@ ���۴^��������I.ho�	3b���,�h����O��Z	~2����OJYL�o����d�@` ]�~u<�X�%7�,�t��* %�!._�y?K4[�*}���� :O��e.�CM�jf��]��I�b\��z�������d~e��FW�R\Oҕ��d���=Dz��U;ˢ�����˯�kϐ�,����0�Ƽ��\Z�ʾ�D�1�e�<��Ҋ;R���at/��v��D���y�r�����#�U?�����P�I^�b��^ܩ��Қ�����{�y.�^r��{�y��}�]�{d��~���@�i^���/c֞7����_'Q_�*x���~/΍��7���6�+�~�_N�M���-�+���|E|��@�ݸ���n�>y�{�'U���Ǽ���v���A�o�õ�  
H��AWo�x�рY~^t���,���Ɖmq` tM&d���EWo%��!l��=�Ŗ��4�HYC ,g+w��:�g�r� %��q7f�!_6;��1��}-��Z��/�L�e>�=���J0�! �@iT��Q��� $�>ϴQB럯)�옌�"��d 3C���"�V%�.C�`4I� ��.��A�+&;�!I���L���whd���ќ�b#b Ό@ ���ɼPn���?;��QL@D�s�y��\��u�U��i���e �OWJ��Esb�dڹ�OE�]�x��#Em������Z��K�e�HET�YV�h+h"���""�ˠ�uW5�*(��a���R�`T39%�[nk�S�\00\�BN0�_/�B��6P�
飦�\����Ιq�<�cZ�FR@0@�U��b���&�U�TZ��\���;�V9�S����*�F�qs�58�EQ)��K2�#fj�kjV�Ėͦҋb�4��RkE6�`�e�ȱ��I��F��4LX�V(Ռ��cz���.!ch�V�L�Qb5m�h�CbmCd�d+b�iTب�"�&�L���Znmj��E-Z-lcV��b�UͫnEm�Qm֍X��6�յm
؎2��-�q�N5%p�%�)_�ĉ��_��Q�pq���Jt�H�s��\j��r�V�*\dN1Q9�!6T�pr���6�\i	΄9�S�h@�LlP��]t�8ԭ��8slD�3�6kL\�0�?�楈��)+K;-*�j*�`���J�&&I,6����w�1ӽSz�8��ʕ���y���+��B�!ͬ��ˊ���sQg{�Ӑ쐘M�$�Ac"����"��UG�o'9�[SZrm�&�c�h��b�� ���:YQN[x�u�NKex�,����L��NH�6-r�\e�[��l�vG,��[R���w��a�޳H�r��bv�7Mvk��	[m%���fU�$��d�6J�g)Qً���ײ���W=��AZ=��I	!BAclF��"�*#2r�-��h̗�R�"D^�fa�x���F�V�&�lI��ڦ��l)�Sb�"� ���3Ȓ.Tv���+��5�K��w�}���ݶ���I8{$�y�۳���$�̙�\'@`*�34?��O�q��:�B����q�5б��5�����%I��-���k-[���Ҥ�gȣ�����,�	$-:�_�z���{� �ǧ(�;����y_�ݔ������: ��2�!3�ϻ���|�A߹��!��;�.��Z�k�q�.�=�P/���O�[�[��+������^�c��K������{rh�����.Y�ۣ%�j������':�o��{�y���ӯW>%��v�8�Sjm(q�E����Sd�U.4��6m���l�ڋj�h�lcM�(�T��cb��5��6��kQWTl%lR�i��*��iE[� #�s��߾��;x;�zsP�� �u�[���W�=�3pq�D*
$�I�g�r�d,ַh+��ZI&R��\4�0�pԈ�����#*�kJ�!���$�%7�}���GII�*��N����g�1�Q�QJ�� �P�N&6x�<����LI�W�-�>�������w��yl�33(�PYPL��j]%��j�t��Q�4 Q��×�5o�[����?!�_��M�	�ry�����z) �L77�--hIUh�A?��3��`\<�h%b��M$���������)�;�ش������=(u��N[��Ѝ\�>B�I5	�?��M�%BJ�ٽO�F�ҟ�&��F�JnY.O5
��R����?O-���)�/SJ��TJ!W����"�%�6o�"�Y�ڥCB�Lzx�i������x�R*���'a���o��@���;�ku,0����ܽ��ٖ���?6�T��:�:٫7�^m�F���מ�<�
�ߠn5g9���]ZL�}������4 �1 �s?\̷�6�]H�M�0�5��AGA���1لp�".�fM =��=��=@>��5�p�싌B�PTdǼ�@z,��*�2"�&2�K�#��� _ �����@�����M�m����
�Pyޏ���Q�<�}�6b7�KU����|]�=/�����!�})s��U>�~t��MI��"���x��M��Q��0U�m�S���D�U�0J�Tѥ���58��<唯���Lo��̲nԶJ#��Mf�\"�ZѨ�f���:(��I4� �1  c lD��T�>&����7���s�-�
�'2v��;�".0���%�_Ê�%�Q���lh��D0D˳#�)��y���f=7($s+�l�3U��m<��x�;������\9�-=����� ��-��d���)�`#�G��0��u;��W*&v�m�uvw�m{U���jJ�QT[lj�c	TV�j�l%i-��ݘ9� �H�� �C��bB6#DXbP-E(+b��dR������r�f(	"!��I�Y���J}�\	�m��-k�h6��5V�й�TW6u�ӻZ�v�˗M9ֹv�\��R���Q;�9�\��@Hdd�D�Fa�� �A�ѷEwn�tιw5��wv���wwe9˶�t�R;���ٵ��:��GN��:wn��λ�v�s�p3�K�ݲ�Eu�\�뺄���1�Q�W!��)j�Q#�.|;�ۋ��P\̣��eL��B?.��p�B�m9)�ʇ8�:�c�)����sÒEz�Ȁu�+��P�+�!�����G8��g\��z�{�R�G����!:�K�&,c�@�k��p޹^9*9�fp���W�xavf���Eu��î.�q�sB9�"-�p�G����
��!6*�AE��H�1l5ɻ�8)�S��w�W$���g�(j6�ۑ#lp3�fw�M:�U�{!��k�(����\�d�c�H�u���܉�3���mEN��"q�:��ǳ*W+Q��]ڥa�Ec�v��:�f㛙�
�Aj��H��Sw���u��0T.��k�����j�f�K��ӻk����-f���j6��Z����Rki7o���u��z���<��L���q�O�i���;���wk�/�����y����q4��vU?����?>���n����~_���?3� ��n�Q�/}礼�'�J������n�y�/��';��i�%?��g�/�2K���:\��Z����� �  '��ð���ݚ@���Y��o��v}�~Yr��_^Ϲ?�ή�)���\�P��`�۟�����3d��t�OS���һT�Ī���z�P�����p���ʑ�N�n׹��U�TT��r�F�����5L@��Iu;kX�Z����۩��E��V����_b׷Ǥ�t�=�NB*l2����Щw��)a�LwzlH���յ���'��)[T	v�Ǭ�(��6�V�ûm�p`�X��A:xzAt� ��1�������Ó�b������Н�p�0��� 3w�!��� q�������񙇮���s��w�|�F�|��L�c� �p��3�ӣ�BC�G6�h�#h����J�jZSO�
kN�dʥ\��0���?�\� �lb�Z� �Uh5��Yf�Y���g�y"9�s�U��������>���:�+Z�j��-��j5ۻ����h�MF��"6)3��YXdP��Q�3�8_�|ϳ�������s�_?�{����OW�>���@m�-�?��=fwe��������#�ii� dp8}�<7%`h�'L�ۣ���N�e��i��4� �Mo�*���M��(q��Dm@ڡ�J�C��m[[M�1S��"�m$8�T�)��q��mGӧ֪���8C�A�&h��n�4��������*
���|ޛ`��g/;�����8v�=�`؄ 1 � 8�auI$n��O+�H�i]V������8��\�cQ��.�3�Z��$)Ow���|�Y���&[:2�xˉ�&�Y�$w6���7)K~���z�'�c#��b��}S9�8��Y?O�z_:Eې6��'&����#M"=S
Y��w��(���<��g_�]�}5k��^�K�b�k�i�+	��豆�U�}y9e�̕:L�'<��X�'�:�J�j�ǵ�7Y���ll��A�Q�m�҆� �H�H  ]zEc���2�纬�\NN��n��%�>�笗�u)�PmO%�K]S��_$���u'�]o8'6|vOݷ	��#���ǖ�'_QN|�IKjw^����P�\�pJ@���\���-�3&����b�b��>S�S ����*8g��`����^ڴ��:�����xP(�ZIiUL)��5��J�m�]�FP�MV�[l��[A�8��yy;m4��kYoM�[�*V�JZ���~�}��Q8������ԇ��6�b�ߙO��_��N3���'��=���|Oe��Q��ìo,_�~�m�����<��'�R�Ha8��B6�j�c-b  צ�m�|��x�   ��!U�!%a���s!�0 $AKiy�{��r���q�=v>ݯ������a�i�w=�'�=��S(E��1U/���:�4��n�|�r����Nz+*��;D����s�Jqէ��M�bG$�#�w2�랼d��9�2��	��F�M�l�1�,�3	=R�6e�G��XqdW*պ��0�=����5|葍{
%x$DMrc��Z-�23.�C��v�\���w�3��;V׹��kֻ��@BQ`E @0�!t�n8asyN���y|�8X]B��|T8�.��T�G��o+����d` r��G�Ԑ��Yr%cc��O4q�'���D您OD䗷`�I��aJ32�u��3�.V�hYs�2l�LA$i�çڴ��]| "A?�Z�e�Hj���e�<���a�`�V�5l�.�n&�-�k_J���
�+qlUDI��Ν�ʔ�SkӭcmX�ȣ���'��[��5}oy�ޫc�^�;Y�r�S��O�v��m��]O���M���������B�s0!ce�lȏ���;����C��{I]Q!�55Z��ʂ�'#���t{~B��mI�}���+�&�j���w%qՅ6��G�b	LǑ@������щ.%��/��bT݌w�c�=��9��>Wu��ʚ��_
4�h\���u$+���6!�(Ǝo�P��Phm��Av�9)O�3��Wz�^A���C6<�v,+A�,�+EY$���ϗ1l	��@�+&��
)�|�Ndb����R��F��R-���g̤z4l?�!Z ��wl�`�Do�ǒ��n����q��_�yk�U�u
᛿ۖ2�?Z�p�>D�0X^0��"�1�p�!�&�v<�,�z������%J9x�d�0t]r5
B }T���e�^K�<f��hY5bl��i�U3R62��l��k��wW�Ž�1�]��ͤ�Hۡ������l�>-�c#b6M��j�jMڼV�m�TQ%���@%gD�1c�`7�n@l:/3���������UWO��8�U����e�����x޿�D1�3�L�HV�,X8���Yh���[���٢���ZLUL������w�DPRd�f6��w`�ndi2&�f/�s���� ���cm�[�b�,�Xo�]�W
a��q~�q�S���H�K�s7����衍���t�o�'tٲi�ѹ��	�Y�+u��f�Fif�.$�&R�\�t�ժ�K�|jfBa�^�Ջ}�{��d%t�68-�GEA���3�y+0���"Bk9ls�UE��"����F��B_T%��q��}p�&g�Nj7W�3�mΨ^D|�p��W$�M���Ee��r$/�-fT]��-dBC;�w9n^�8.��J�wZ%C�8���4�p���nX�m��k7�`��,#�7p���C����G#�~9�������:�v���eוǖ�	(��� H+3��w�j=�n�&��8��Q[�]���6���"�HL�q�9]�ʖ����o&�#�(*��*�w��촦��ř��� �H�y�o�5����8Q@A�8m����_�|݆���w�~����e?�m���7>������=~ˮ���c�g|9_c���5��D.7(c���+[�_��o+�/��%��_����U]V�"�	ND:TU�IT�:���##��b��UDrZ�JYK�����hf(7�x��#�*�KS��%N^�Qn��_�DƉX+��x$q�� ��\� ��!c����k�F���S α���h8�nUٍɻ��%#t������V����o�9� �Ӯ��B�s�$�9\����T��Tz�6�4bRK�N�U�Y�dM�\��(�Uo�r�3aZ{�uʵ���\��:�&���W��9�o0�wc&W*�|o��fr��y�T:��ί-�T\E����U��h^j|FmI�NLD01l3e�.L��!�lӺ�x�p��R$��*���x������Y��y��IztJV�z}�q�Rbu9���u�Ƕ�%�ꃤ�+�+C���֓�8��匮�,�7CRd,�kP@��!L�ar�<έ�Y��Kpƛ�{m��ܐM{_˫k%�)C�e%�d!*B$4���ox��Z1����n�p#�Ѵ�ɴ��[J��t���h�b�wK@�1�K�T*,U@8�+��s�I�9��}�]�q�F���]'���=��_5��鿷��y���_�W��������������v����� �4 �"_�h�v�����2��LD�M%IH��A!b(�i�e2D�fY2ř,�� � @��q�O��5ޣ;�r������`o�Փr�RoJ�԰�	� �D0�|,t�L�Ef��W���r5��hW^>�G��KGd���S���ѩ�wM�^��!U>3�-5y1���3�]Dˊ�^2�d�j���� ;@r�+:�r#4�*1X6�I-��8�<��(&����z�����+Ӧli|�Wȱ6�S&�Őu��-��j��O�5�$H9{��Bm�KT�Fst��i_��P|�-A�S�D�	��yI��[��0����q�sF�9�:K?�W�z'�d����r��C�>�~��oW�N;�Jo���@u��u՝4ƞ<�yA �ȇ\1-��l�-�΁vQ��2�v�<-.�pڸ*��6��^ML�J��T�Q$%T`��Q�����j]w��;/��C�~{���8_;}�?���ԉ��l�W��g=_������G���rMp ���}��h��o���С�����s6�C�Sܜ��I��=KT2�9wArwE�K0���x7W�����5�H����jT�0B� ��ұh�Aய4sdW8#�9k�;�L�Irh6WFNP��n��.��U^ҙ��/Q�����ׅ%&��t�K�9I8�G
�"�h�.��.�α��R�H�ixVB%�N��Ρ��;��J�n����DR�wd�F*O ��S	*+7W+�\�P��$b3Z���+#E ��BUC�A�增����D���F�wT�"y�nWjp�3'y�E	���j�FQ2ĉ%j&wQb'����U&�D�'��#�$��:�$A�]T<"�+�;�WIz
A�=	%v4�p�T!�y�7��*n�F=��T�����J��n�
���'��L��ew�ITU<��)̭�)��D�0���Bû���ա�X�^�bR4�C8&����7��ùQ^�d)��$�7��(�hK�*4���8;����XU9��:<*K���#��D�uH���s)H��b"`�Cj��Uu7G�wF duI.�r�t�D6;�4L$�˱S�w0��fM�V]"f�j���y��"�D��;-^�2�[�j�[�!�"!�³E�w4X���*��F�M(����{�T��"�%�����h��5JOxj�=�pMFeP�'!�,�v���HW448c
vJ��AT���.p!D]�x�"Tz:����0N���QկpT��Jiy�n�7�[-Jޮ�
	��.�xS�D��j�i'��CvX�y���=�B�"��j��w"C��<J�2%!���V-TWI������^%$Ќ��#�SEVt�t��ttZk�XC���a0�0rF�,T��Eޔ�h�p�n跈$;�J�"(*����H栉/PL�^��TIaVZV�os�:#$�	�
�F���5f��,otf�g!W�Ky�$R��*Q�t�53t�es�0��l�tG0�m3AI,��ƨf�qT�5y���B���M���BoJ�W7grW��j���9<��8�ء�R����nU��W�	Q{�J8���^]C�I%�.�n�tQP�$QNP��*b�#ѹJ�̳���+�+GCAF���U,�J�ƧF�zi��"�Mf3�:�#)���"��b����L-5�$���IXz8qJs�/G4/,�L��wf��P���]!��-z4Gi�'�L̈h�K(e'E4��J�cYg(���S�E�Ѫ��p�Β��p��s�zwuX�����P��3�\�]�j��\�R��"+A#�I�鍈�%�n�4�$:ZUJ��/�G%`d���]�̉��(̕.�A� =�Xz��îT��#���6i�#r���������b�F��ܱm%cT[Qh�b�Z6���c,Z6��Ƭ�RE��fH�	h���Q�(�[ch�ETljMh�mh��+EEbJ���j-��-��ƢѪ��QY*űL�6�c�,Ecb�h�ъ-�ԗn8�ڑ�-��k���rޜ븸=MU� D�K��cL���fsK��en���U�Z���l]�E4!�+LtL�ٽ�I�#��.������Α��<��IK*�XVw[�����/xe�{��;r�j�nMƷ;�H��(r��/���ǡ6Վ�Z��u7�Bً�m����2졾2��Q��L�S5}!����p�$·S,�,�U�F�ֈ�I�Ϯ��{�e�%xg��K�n9MeOƩA|o�^V������G�ݪ���oK���f|fxB��[�^_6�Qd��9NdefgZܡ�m���+�Z�gL���pk��]�ЎJ_���&���&��(��]m���[0��^#WM�)�T�֢�W+�*
6I��1 �c�Z���(��J/_��]�Ó��?�����������~��p|Wg�{~��r:�C��4�nMb*j(��("�R�;���z�.��D�эn�d�Pi�����lnVm�j��6��Ø�?p�4�������������V�7��2�cN����P�|��D�o�o��MkOS����ط��lk�ʔe�^tr<��H�������Ȭ�JI__��ӕk��hB��_L2�r�ga����5
f�����`�����1�5��%�*��/<�Fu"��F)��qg�5�+�r��ӓ|��;�Se�4۲+-�#{�֊0Ʒ����?w�٧�����rs�f�>	L�6�����s���xpߊ���xߖ�P�M?��'E`�k��Ş�\؛y�������[����]#\�r� �b1�_��a�����Y͡}'����o�E��}���CU���η���|��h��=�� �m Av�24PJ7���ݯ�=��E����T��OҼ�h�p+$Ջ���(�
�Zc�q���yXY|\;h�2=��	qM@A91�)��kk��wiz���b��;��r�QcA���|�����?�����_���xC���6��[��CS�_��������G�6�;��{~����~�.���k��F��=^J����c�XA��,UB1���n�gx�>���ۯߏ����:������4 㰰�J����-�v��%�4�Gx����	���^�j�nsE�cBCb��*�o�?��p�r���G�������#��Gu�;�;L��S��?o�����|]^���۞��}/u�{/�]�Q�7md	:�F�
P���5�U����y�A|�qt�.�CU<NB�{�&@d�H�]eSa��fk�-��b �Ͼ���z�&����K�s���u���o;ƕ=����zݎk�tY��;|�}���1o���s��H*� �`��-�Z�̈́ �t��V$��n�V繍Z�ڮ,��PfLJ�� "`��yv�+�b�2Eߝ�{�-�������w���y'~������\g��zxR�_{�{굔����WQ����Ulv��f� c ��C@v@�z��k����"HoTv@fc&���c��5S�H���C>�2�_��Qs�o�
�������m"y!a�0[!����}�׸
<���V;o�S�N2�?p A���]ë�R
j�D�������b�.,cS�T��'�����r�d
ۙ�#=\��\��R�O��J ���V��́�ه�K�ww=I�C��\�C�7�p|��=s)�߭��|X�3�a\�O����c��_�����Y�Aq��H�$���W0���NL���Ϋ�I��,c�,{�vC��Jm����l����@��Zޗ^�y3�n�}�G8��a����Z�y2~(���Rm����W��y�ug�����Rl��B�d��?���!�c��m���3��sv���sf�9��ia�n���f���k_����S�}wo&����1{7iF]7��C�� 洿���׏�C:G*�0�Gߝ��|oo�}�4�ZM��l�6�;�j�<'3Ms����O����y���<�n���f���n�N�l6��v�y�/5�y���<����v�]%�9_��o^�ωid���-��9��n\Ke�ޟsA���7��v�\�i��=B<���n��!;��7y����p���!�~�����C��z��2^[��k���ѡ����L�O%��ç�}m�R�o�4�ξ\�	<�y���_^���6�'���寉)@��������7n�[g��w��=?�}�='#"-��ɚ���o�g���}7ɂpe�,{=��̇�B�WI��d�Í�� <��ֆ�!S���I9w���H8DX�Y��ih|���߻����z��|���ܬs�n|H�!���T!!>!�B�.���L�D��m�*8��$Wչl��rbI�/װ��늰U6�&��*�s��vx�C�X�Srif��}���s�m�M��i9�}T�vSHG��/$J��]۲+��Ӟ^�w�q4�f7�ܯמ�lNRNkx[Fp���^��7BB�(����_Jr�]���/��s-��{��p��Q����r\�z������=xs���:Q>��ԗm��sw^��}n��0ؾ�{���iH)n�g{�S������O9j����ۗ�6�<������%V���<��&�Z�R�qӗ�r�w�[�wl��7]�O��N�3ɐW�'Ok�|�� ����w����>���.S�q������,��%�ig/E�Ѷ*��Wͷ9Ѫ�+BTZD	�̌2��U������J�Tji+*�Ed��s�<UZe)=}q�~7����:խ<�h�M����������KK�;��-k,k3,�����U��ld��T�E�s9e?��5�uu6�U���2lf6Y�f6���'u8�je @$F�US!P�t�����ɘcP��S�,����������������Y.f�:8��7��χ�����z-0�x4�M4�X$�6����-��^ˡX�LJ�*'i�~N;
�kG�4��{���t���%��2,�y����9oy�s=��i�Q��a
�A��$Hc1�������!���"T$B�%�Gu�q����eH�A1�����%�@�I@$FGn�e��g��C��L�A���0�0��C�k�nI2�H��v���޹����xBdMڧ,�b)%R�'k���E\�[O;��d� ����2umt�q �M���v�����ŧ^�m����$!㲛��Η���cO�۶�m�8/�%؛�ϗ����/����!v/� ���
H�!�"�݊!�6��K�zo5������������7����w��?�JǤ��(�#��B|��՗M������=���]��v�x��������?���k#��^쭌I>DI�����o�No��w;t����m�ۥD��>�YXUhF̏�7�&����k������_�����5G2���Ǭ��o��8��W#�-S�G��>g��Y����{�g20�aU��9Y���YseD�/���U��e[Z�J��ŧK�D�6*�IY�����~�oz�M��e�q��������(��	k�M�[��^��q��i��4Y͂o������e���tW�#.��B�Y�h�S�ivSÕ����G�m1��4ZM��&�:�i�����ghlV�n-�-|=��4�$lm~#gh1I&>�h�lp�Qƥ�
���5֍�����&�4�K�8�jc��z� Al]ʎn :Qn�c\,�`���* �8�E���m�魻�OY��Eqń� )(���W���@��
bS�Þ�/�ꢙO��>��2ET�4�$dD�}8Kq1�V���U�]5Y\�J�.<`i"�����a�>p��G:��eny`&��Z�A��t5eoI8?��q:��:}��G��������o�!�L^����F��A4��ц�~��\��k�9b�!�����i{���a�\z?$���s�O�z�_z���y'��m����� �_��wG{��'�V9�;<y4dD�a@��%>�"Fǭ�:�e��0x�+ՏR��ҝCx�b�`�b��b@P���m�C��1�q�s|o��: +��GM<��q�<0��l�����پ�	��rAP50Xv���� ҹ��p>/Y��f_٣��M������@r�E�=E.ci��]>�1)"2����7�N��wn���G$��k�d~6��� 0�2����<O�����f>d`�h��in��D�X9X&�E�P���	�r�._���K�û��2����e���(125�����_�
k�?�z�F��+��L:�f���?7�o��)�/�ܷ=���"�����jH���Ӛ{�E������Ҟ�&�i]���8r����\�����~�����e�ξ��d	e��Aݿ��š����1�{ �u�}��)��V�#�)�����ӻ;��������UQU�`!i�?�sw���E�m��-��6��j�&`ڙQE�M�^5\����F�r�jKb�A6M�sWwG �#L�7r�:Rv��3��˥j�mA�Ed��Q�H���جX�6��"�F3,cF$���e��3�3ﾐC��Q�,c�2m�J�Y�V�֒�E�F����fk�b^Dr
	-/7����L#��7 0$l�ÜM��rffs�d'���	c�H���W�ʝ
�-����.�Km��N{��H|����HJ����X-�ݲC�iXq���F��YJ��Mn6lv�Mܪ⣚�r�����x�2��fKl�o����fPEAz�;S�^�+��t6[x8�c&x吶dH+"��`ɕ*x��wW4;�<����L3�Рx���"�q�����ݎrK%;�wrPn�e��
ws��v��.��I��U���1����x��"�b�E�7p�6w]��]s���F����]9Gu��˭s�;���]�I�a�FF8� <z=�s]:wvr��t�ݸ]6�r�;�;���r��ͼ�����'.�I���8�Wqt�s�""��r乻����cwt����:�]*�BAc DX�$�$��둜�˕r!�t��ӧ�7WL.���]9ۍ���g���ߜ�r�*��.�����D�h�"?���ׯ��9𠾏RVO�!SnhJ�eZER�l��ie�q�e��
��b1	m����։�I&-IX�:R	,��I�.6l��p�� ܷ�rt�EY�l-��T�V�����W ��I��ZD\�Uk�* ƣq���K#e�l�m�Ī����hfff��w��:�:�m����E��y��`���ht6
a	D$�HJ����j	%���Ҁ�+�M��"�"�L"f5�kl�����|T���>;��.�Q����$j��S��!��ۼ��vnڪ�ڰ���A0A�YI�+$�H@��ffFH���p��B�IP���+�eKݮ0��9.��_^7w���%�E]~RW�'�6.G#��5��a�.@��K�b�Y�*Es&͢�QMs���sʋ��$�ؐ�֜K+/�&O�_o	�G"�������)�}�(���a��58�"#�vdپm���?�p>Կ)�f��6�rL?)|��LN\�m���[�_<���2�wQ�/��sq�s�r{�� 8q��<���-=���{���f�L��d0�r���<�棁�����'�������ɞԴ�u ����wo;OS�R|{��o�}{r9�y����{'�=��Td�����ٜ�i�	�5&{L<J"5&d�2����'�˻���۸i���>��W��`{�O���g��
��y�<a��E�{|頚&ЂT����ˇ����v{�L�k�s���\��>~�3B��q���"��e��H̸4A���\>t�){790�[���<C��!�޳s"+�`����x�����L��̴\/�d�!��8W)īI��E�3;0��v�I����\��1 �)��+�e�@�r|�W���+g�m�ru���n*�>��!Ɂ3<~neω��i�%���s�܀ �d�`��$��vdGeID�0�^���v��]�o:�)��
���9�n�&&# ܙq{��HW�����{��+�����B��� ���	�p��.{vd�|'���â� ]���d��O?Bg�	���;ך͆8 1�=���fdO#3�\�F��͆��>[���;��s�nX���	!S��y�L��˞_=hh.8��S)��pN����p���NN$ݛ�7n�J2m�B�0u�&����ܒaWy�N ���g���8���=�|�O$]{3Q�t��a��n3ڔ��'��P�=C�t�|B�|gxY�^�#��1�;x9s��̉^��s$Xt�ԩ�9f^L�q!Ďb�E>�\���ϗN'��'<Wϟy�����3]ܙ�MI��"o�.>�~P/;��zq���㜐QG�1�U���$�d��cH��,$Q���ps���T�}�0��i����0�
dF�h\,&r�ul6plCi
#�Jf�i�|��9�l��T\ vf�3�u�s�T.!Ʉ,��N��h���20�Z�D���7�[�<�j.=��9�P�d�1$�p��sC�_Z9�v�0w8�E<�@0Pøv��T��0�p ����IF��W����۴�3���|��I�t
����̟��}�[��&�����.�LW��٢��%�_�LU��`JM�����ˁ��C�}'3�Xw�L�ߎ���6(�{sJO���s����#{�I���V6�O���B�TB �FI*�a+n��� Ԝ��	��E��\k�w.ve���=����
��ɲE� Tx:�!
B�X�S*�������uwsk�t�nn�H�D�����o����zp<p�Ď*1��ы�����oOg���������x��w�f�}^I��PV��m����xcDbF�	.����:���w�mz-�ֹ��\ܴQcI�K�Fʳh�R����Ŧj̱�l0}�޺U���� :��@`�m	�U�1(@�ˤ������?��K�m���z�s幍�F�����-E«���1���Q*"��B*g5,;܌��z� ��}J�a����� �Pc�g�-��v����[M��*J6 ���lj �H��"O_w����� ��F�Ha�EX����ӽǺ�����ދ�F���Y��`a՘�/��O�d�I��2D�\+���g)\|EG���������.�~O/����s�d�d_�w���O��#;�a���d����*,&�؟z�m�e"n>/iXꏑ�u�O������ߟ�|/����?[��L���{,��{��v���y�z'�i�pd��;�s�+�k���X��nk��~��'���U�4��@{����'��?�U�����a�3����.Oܥ���o�����S��WW�w�=I,p�yV����v\ݦ�S���/sa.��GG�;F�7���f���S��}�ߴ��
�����l��ʉ�F+M���}�g�:��ʕ�p\���
p`��s�n�Z��s��T5���{�.��䚇Ok�L�q�+C>nW2ζb>$�W��t�j~u-����<4]F��5�CL���1���~�G�-�dg��y=���7�h0�k_|�����g�����S�o>ί;��{G���qki:]���ʽ�;O7���i�����>����ȕ��#��8�Y����e��79����>�G#��c����?�οoѝ���4[=�ힿ���N�J�n D Ts��>W v����x]0����o��3?����m36Wē�����?�������n��C#���E�^4������=��o;h������S����:7u���I�����k�ɿ�}�t����p~9�
��x���3��?S�� ��?�rr���>�ЫP���+������U����t�����֟5�9%�8�kg��5t�o�]��K��/�{L�zY1�����z����$�] �E�D����*����F�ߢ����i�WA�����Ҷ�e[')�7�[�$�0�z-�����먿jM��#𰜓�ZM���HHO�-�ұ��S��)��ӱa�|O�{�/��ǷR.F��;?��8! ��d�׺?��s���L,���hM��a�.���ƈ�������4އz#�e7fl���u����@������ޏ[gk�J���n��]%���=�}_�a����~�_�������rTR�3<٨�.H�BFl��ʊ?ңA�?���.����Y>{F������?������_'����tّ�O���}�u����O���J��0�*I�g!�x��mUP�'��g���Hf73��~A��G���Hжb��T3.�E	/�/C���WNv^�sJV��C�.�
�J�a���9a��=9�6G>��wI�ԓ�OK�a�ge��|��짞@]��ԫ�����֧�������'d��|>�M[��m�1��O����G���&4�0X�&HZe֊�J�ŕ}R�n�m���40�fE��ox����=2p�GO�tMt绁��e�"i&�h�_��sj�yIw�_�����?���G����.�U�	q?j���.@
@���g�ޟ90��b�+�\=O��nH��! ��y��| �;�?��� ��>��Z�l9f�5'm���D�����y)�65"�2(���)s�yӸ1zq�P��+���}u���|}��#+!F!f��\�X����OAб2"|w�C` �#:�ۭ��ĦK�>6�9�֜�*�nCq�v<���F�7�����6��u�|{w(b���<o�	���h1a�+����x^\�i��z|�e�2����7�<ҋ�u�����/	tbx�aA|0�m�w�9hA�(r����Mg(K2�8zsE���=`�/U�*�����m閦���;@(w��V
@$d@v_&ٜ7\%.���Q�uR1L`!�x�z�xGLu:_�{��7�����u_��ǧ�W�z��~���!�������'���8����<q�F�z�+�����,�����|�����E��>݇�ߙc��?���|^���?�ih���(�~��`�~?�?�=��_o(�}�:��]����a��9�}���ׯT����vG�o;��\����D��Z�m�6������͐_/����+��蟹�Y��&��f��Y��x>/��ya>bo�.x�:n��'����;������_���}�к���G7���W7�����yv����[�o�{��?7����-^�[���>W�8��[�I��u%]S�l�SS�П�s����2�����١�|o�ع}}>E����<lOO���P��cF��8"<�z^@��&�f��2/�_�>O�B�Z|�,���N�W0�#�]oCBV�A|v{6=�3N:�4T�����$&�JvG���p�n��#vȿ����� 鴟bw�����]�$���^�*ӥRȿ���\MZ��%��Z~m���Q����������C_G"vu]n-�^�:�݌�������k��x7�	OU{'��ݾg�+�����W�r�g�����aI�"�j-Y��Z�&4r%;�.�Jӵ��|rq�[�����{G.�U5F%����D�t"�J���tx�4Y�S̩���K>�U}y;MF�[��YI��n��1-1J���>�.ǽ�+)�>��r$a�k/el1�i�WƟ�el��39��D���[�kd@;�����̌q�bg�Gi)C�G)Vy~�Zn�be�9۸J�����~��]�h���=B���Օ��=�΋j�3���V�R�j͜�����\!���~r絧v\̾�ONk��V˅���G���̚�+��{�_�?��}�o��s���y=g�=o!ӹ�ߓ���s�_pڦ��;if~�y�����C>�Ȇ��T͍�Ȁ����������	D����r���{gt��<=���A  ���QkZ�x��7*�.%
���\��P���}�J@��Χ���WtN���8�~���L��o���=Gr��m�fW2�����9?dX���J#��4���_��"{�Nj?B;;����q�RZk����(���"�;�����`�"D[�M9Ӏ�ksR�R��c�Ї���v6!����H�F�8�#T��j���sz�3��DL�P�ѐ}V�,=��1�>����!�Lja#���n�(��n���a�Ϝb�#6:u(�Hf[�H�5��gMFT����%�fL`�Nb�Z�6#Xƴ�5�Z^C���¡5Cl�)�>8�a���:Jq�'PűVY�(�,Y�'#r,X���v��^,K�����*��\�OM�H����54��u��cߑ<�_�9H�.Mf/����b�L �?a�N>�[�M"(?)���T�(^j��_澖^R�m[/���ǜ^�J_��N�ta�sP.3R���[k^�3�Huf�右�!�>� �F+��1�Jo�o����g�!��R������{)p%��~m�)«��JR*��)>��R�-���� �l�U�0]����'ҿ�k[07�tGs^>�Om���ι�2BW�a��Z���G����\ V@'�8;)����+��	$$�� 8M���>b�(�`�FK~���6:���� @���R�e�{%�.;���R+�����������p�!<7�wQ�˙\�I�F���d��f�6C	�����l'f@ڃ)Z������ڷ�>���.�)��\�r9�q�^��y��hQ'��I���xݻ�*���I*����C�U��ƀ���a�9�s��c�`I���/ϗC���?Ϳ��S�.��U�m���`4j�Y�MZ��a_����?R/�J��W/^b�J]�pJ�]���|m^��m�eЌ�0DL M��oe��Q\�W"�4��W�vG����l�iWUXF2�����}9������d��?����v���Z~�-�/a����B�9�ؿq�yȳ�ݘ�X��ZhX;z)�%�)>�.�2�jnț6�D]r8�UUU�Z,�&X�L�T�x 1��^�\+���S����%.�y����P�� ĺtG�������Ȅ�H���Ւ���ZS+iܡey~c��t&��@��L��n�3v��m�/�}9���ϸ9�f��'|�r�(�j�����Q�Pz�$K�.~	_��.�l�X������� 81^}y¡�
���+��B(^ԥ�䧼������'���.˓���*~��uY�ZwA� 0߰Oω�s�)�H�cQdѵ~#k}�v��A�ʺ�g�TOTz_�%� �(:��^�$�7��\�B$d�!ăW��#&#;�II&D$���ۮz�`a���l��٭�5��G��R���_�����H�ỡ����(�p���wɞ���w����������lp~��o��~l��|�^��6��W��O:����Iq��%R���T���1�$`�n��ю=��IJP���6�a ATCgt�N���_�����֩bߒ���ؕ>P�����S�rq*�M�j�
Q�Ӟ��lw㌾�����eu5��T���nHGP�K�~�:8c���K�|Bw�mU���(��O�?g4�����M��+�y�/;x�����>�1�R�\�O`(t@���j��s¸G�7�Ӧ2�yW��'�x��8�2����*������^0�/S�I^�Ҟ���H���M��ݣ3����U֖�����x�G�N��D�iO9_wð�ϭ����C͢�
<�	:�Q��ާ�|��u�OX���(�p�3�},ƲH��!�I�A�	��H��.v?#��׬{Ce����66�P�A��0	{v�>�&�UL�*���P���1�m)�B6.�	��`p2@��W�|^yS#�z�~Ej�.����P
0\��Z��C	��y��������>@u�5�ck6]��%B��#���y�r�.o{������Qcc[���M�����(,��;Qws'km�WW$�I�3p�7+�W.]�Q�\�F6ɤ�5wunN��:K��q��L$ILM$T�ׯ��q���^�:]룣�m��.}d����N�W�t���/��v���qBp<�[����X�fƶ���x�.�>1����x�r���M��jR�5������Uץ�{!����
=��/��t{*�ye|м�������.�+įyJ|?�^�����*"#�|�B9������������~�����Ղإ�T�*�CkL6���C/�u�
5HA~\���T���4��?�<+�d�hm;	y�� 
���%�?f�R��w��|����}h�G/�˼H�/�>��ҽ[M�g��i]��"��8rH@��a$%��.p�z���/n�����s���i�\}�ƺ/��G������tB�+�U�8��rN)�XQ�ӵ}�����S�/g���G���<qUy·�Y�tLF�OF�(�b @�]p�a2��}�����Sa��b��~���g����c�,/���S�����J;�W��f�q;O���ʚ�&�eb�i�ْ�n{�'V��.�Qܥ�ܧ5[�1�M ���,�\��/iQ�/{�lp�U�-��:�	�Ug����E�YB��e¥s���8z���R�����ܽ_\�(x�?�Sق�?F/V�%?t�(�%�q�+�Wp8�<���
=��๼�ܺ/N�緉:>V�QR��u�Y����\�y��`
�q��1��g�C��i!�\�M}&����LͰD����t{5��t�^h8�C`c��7qU�}�U�X\N���}�q��s��0DQpPGXi�<M��f���������O�S�Y���PƓ�g�W��{���hN��]�<�̪q�(O����:^x�]�t���m�{�8�V�4x�J����/�$�pW���ŝ�)��	�f!vdhH��?����2H��d�G��0�{��f�V��xK��*1i�X5$��K%"��w���أ��a�I�R�]Ǟ����vG���Q��Ww�g��Ljw�<�	��1�`��2�Pal]�BJ��U��cd��z�dY���e۴݊�`^�(d� 9RLk���cRҰ�xR%D�������w� #p���>W4�8�y�®���S[]�z\U�.iN�C��y�B~���z�tܹ��	�Q��C�TDG% �r�f8��G���6R�f����yg�U�����_2<炝ӎ��)���;a���r{l��¨�<*��2�'4m�8B���F�c����E��v��܁Ih8?-�x��ھIm��	��	����z翅WA���k�}��wP�m����~T�h 6ZD*�.��J�E�pٻ'�o	�o�닠�
8}�j���iF�`���'������a����⢹^�U����D�/,6����%�,[�jP���%�������% o!��^�bwL{��j�������n>R�t_[]��R��
>/[�`})A�/���6~l�5Wל�Jk}P�l�����H6wg9yv'Ņ� -b��>����ԣ$<_zS�T��W�E�i�8a� �a,�p�@��/ф�y�g�-���p� d�� K*o`af�rZР�x�g���	Ã�1��=D$���S5T��� �����������Z}������`΅��gV�/�<���\i�,� ��ѽڹ��f�Y��&6qU�^�(����g���"@	 I	��?a��x�A0����
|���x����

#�`�Q���tǔI!r�.��/뭩���)�G����U7�1�M�&�28`p��Z뾥z��`6�[�?�Q���`g� ބ��t^EEduIG�8S�'��_��n���N<frv-)�?<(I�QI� 6bC��$���=B�"uxD��ד?U��0�B�#"��6q!�¾����K<Y��&6�$P�_��۴��ߞRa4m/��������.	�H��5�@�#~�����K!��BS�W����Y4=��솿�x��Pq�B@'�
6��z7�;9��]�&�tp�Q��(�B%������u�1A��n�E�#*`�\ �Mm�s3�Q��'��l�	�20��{���}�BT0�ԡHl�����EB�� 7���u� ���@cC����5����
8�&��+S�'dIO�<�7���W}�kך6��_�[ܵ~�zW����P��w�j"��QD��s8�����?�������;�=�z#}_��w�����?��3��^��E+G�i�|������Y�?����6�����_z�xv�?_��p@p�����wK��X��Yрj����z�=ǲ�j��d�^j9��qi�����Vi��Ǻ)��ս%����W�Z�ix��ﳰ�+����<P���zS�o�M
`$��\vtj��>n+��U['�I v�H~^o�$�������^�Tk ���̀;1�K|6n�W��{��_��A@��o=hq��C��E �d��[�[	�04$�U��,�����Ha,����o�).�Џ���%���x"8`�m���|��	΄]��N��P��&A�l��]��}��I	Xa�����dp@$Y d�!����ޥ�	���m$|x8�����rьCԑ� �F;W8;��O�X�I�����˟����F��?iq��u��	?�|J��:;8�N]�a� ���/rN�#�y+�n�*�A�x�ϗ���.?��IA����!@h�1/$���`]��u�ܢ�@��xlo܏�J���Ro_�,�SG\E|�t���F@?��R�B�E*�B>�?�$/O%>k!+�8]�����>��1!�)��8{����i�,�հ~c>��U�Ӫ�r��>�e�Δ|!�r�5��jhCџN$(p0�!$@��wݕ��[�">z%Gl��,� �r��	ȍ���F#�,ژ�/���'�]$��vf3YZ�e�i��I����c+1��o6G�^DI'N�"�Y[+��}n;�q8�l���H���~���{��������y��g��7��oێ���?FmJ0b0�o���?o3SF�d�QoIG؀��I�i�zJ�8�*�cL�zFp|Mt�#��&T�놽�����I�����R':�<dƌ�vW&��s4IXQ�����6���� �K�D��iv�[F��~�SD�{�cΡ|�<��&{���n|l��0^��؝���܁9E���=����ص�����]0`�{�J3�y/�^s�ӷ��콯Nv���]���e�B,���qG-G��Z3��VV� =޿m,-�B	��Jͼ��( �!"��#ܟ��YKڒ�LҖJ���o�վRm�V+cT��Ɉ������]C��m��lѲlM��g`��o�?O�O�g������)�ru��Mu�UV4��!F��88�
f"b�<�؛��?7���t�y����_llk����|��y���A��Ō#$ada�����{3�UOCv���ŏ��	�q�rI�er��+��ђG煾�������+ ����������ꚿ�B�9��>��8��ܴ甡�L��U�7�SH������Qk8b 
�� ��1���B��~�C�eA?��x�J�g~�{ W����#�Z9����{��M������:*�X�f٨R~J�B�"#$�×;\�9�^��k�})�d]��B��Q�C�������,^��(�1Z��ˌ�\�i��M����Mf�i����p���_E�H�5�Nǎo7u��IL�DF�eC&I%(��&�#Q�A���4���6&RO/4��M6` 
��X�@�Ǟ���K�e.\|�oX���7�==+����ٿ��>��5��V寯��Kд��ٯ`7$���J��b�퀿�  #B�1 "l�J����9����3�$��yң���z�A$��<�Nn�F���͕,�
�	Q,������7ˆa=]��A�I^>~I��s���� 	k �`0 �mG9Hb1��_������y�Ȇ*�H4�f�ӕ�8��*O����C9@�Qg<�+�E0��ih�r�˕�GB��-���q�W�b�(�2�E؋Qi+�l
�`1�2@�"!b� 0b�9�mAT�������bŘ��ˏV�dA�T�<y����"��?LY�"��p�E"�IEH�S�OT��iK*QﰔƟ�|1cDYc�=
��<�YUcT�\����_�~����4�i��VHB@��bD�0������è*2�JfX�~���Ds�"����.�
O@��M���/F��F�+�9,RZr'R�%)����&ʳM�\�����MD��-��MV,;��7�YA�9�vqB$A�����)�b��gV>4�2�Xq��T���M�I��^��j]��n�	lB�IR�ʊb�M���bW��-���{+�f��iR��A&϶�jR�P���*'�!AVu���d�l��2}���X�!zH�.ٱh����.^߫��i��j+�g']>FŮU=�0�}V�ݿ��D���%�,���:d�s���.m�%"sR5J��x�RZR���u�5x�1�3f{xQ�6�S*�X��Y�N�R7*�j$�Ȇ������+�8�	Cw�(��¢��PO��h��b+%�mʮ��r��mF�n�)r�q��N6�B�餬�HF`�G8�J��S&��mv��]���*�k����+,���ʳ5۹5���%�W�͍Q*�x�b�h��6�l*;��y���k��m%Z6�F�sk���m͹�z4��alr�\jC�8��ګa6Emm)��C��Y&Ȳ��.tF���hm"l�©��H)6T�m+h3UVĖ��)�%�Ԇʫb����VҊ��-�J*-�(�B��ډ��U�(l��R	�"-��e�R�U-�'9*��V���q�ʩ��D��M�q�[��-�\���j��(��Zѭ�ۚ��(�5�m��9v��1�Z���RW-�nUx���ѵ�5k�ݭ)k2�cJV1�Ak�9B*K��Q�%����ZM���fj(���i�*DƌH5),FH�VJ�T�F8L�K �)�b��Ţ�1��E�DRF�r�5sW+`����1�1Y�w\hѫb��5�`1C,Q��Tl�0j-깷+nZ*4�$�lljKXb�ٕ˛��ѱ�K��
آ�m��2 k����C����t�O��xܯ7�fq=�����gk4~r������=O��;o��o�|?������~}?k�/��x~�q}�G���q�̻ۛ�~VO��G�SS�~����~�N��l{]s��p������^��_����m_��o~��{���Q�=���-�w��\��x�G���`����ϻ�l�'��:�������P\I$!�Oƻ
���ɪ5�!Lcц�9ٍh�Q�V�e[j��1�bmI�L[b��M��M��5�h�ڴkRV��bѫE�f��P�5&��j���PH����Q��6�UU�DE�	���ƨ�$�h��Q2AR[E&��F�cZ��61d1���6�V�@��F�[6�Ej6�V-�Q��6�kQl-�V��Vж�d��Ȗ�6�m#a&��؆ԕ�-��"T�EmT����"�d6�M�j�ҡ�66-����"�)6��!C`��U�l6��تSbBm@�*�I	�6��l,ʋjؕ�U6��6��!�J�iPڅ �T[6D��Kj(m-���V¦��%[
&�(؊-�Ҋl@�JQ�U[A���	�d���6I6���6Em����Q���-��T��M��i�iJڒ�	mU6&�J�%�6I-��j��Fm���jJ-j����i���ѱQ�A������F�mFQEH�i"3f�4��F��P�E�I%(���h�2U����j�Զ�kf��0�ү��Ԛ�9��4�	W-����?�[W�~.?�}_����GG�߼�>�?��U�u^����ܟ+��~�o�|ޓ��O��u_w����緗��:�#�3]g��0�߳KC�����>��'����?K[�lC�y�����ע�������^����_���������k<�����kQ��x��K�:׻�������t'�t0~o���~�fk���8���l	������gE��=�ŕޭG�n?���n;Oo��ҽ��ŗ��]�k�T�|o�����ۀ�@+ ���z|��(]�66��3F��b" ��)Qh̦E1�(,�X�Ii4P�f%��"��ԩ�(ř4X&�M��L`�1�J�6$�34`J#KbB�Ȧ�C!% ��C4`)$C""Sa$Y���J4`M
H�L�J  ��z+�wt�	
�I���`X�C$���FIHL�Q�0���d�34�cS�e�,�@�"�fCB��Ɉ��Bi��BDɀb
 RHȚ%Ec&�H�FI �����K��� F�K�"Mēe�H�&�L�(&���e22��C# F)$�I2�$�Jd�2"%�@C�d$�a1�X��)"��4��#@&�Hi��B�ƈR�A�4�$�6�ɓ$ČHXȠ"�"�ADa
�Q4B)������bb�#E��h!����L�%
0H)B�1A�4���04�FC24��B(!"�c0Ȥ�,�����R�T#	 $J̚R	M6,���F0�B� �2%E� C�D���cF�4�H&�F1`J$`�2B$�	�If�Ȓ�I��e"XAIP,T	�&DY03JF�eA� ��>������m�N��o����=���jk�j7�#��W�^�Ӿ��~]J}o����_�W#�yٵ̣�k~������$�o���;��ȇE��v���>gG�_�y[~o/��䀈B��ۅ0���۳�z�^��w|��r�_��;^���q;����������]�����26������֯Cʭ����=g����!�Q'f�/���n��{��D�\�I{����>׍G���s���}����}W�O��5"Ա��&��G����_j0HC�=��{˜�'��&ӿ���e���v��!�������r��cM�������f�X�?��fwʝ5�?iQ�.�T&O'dJ^q��$��ʂ�Z圙�W��'|y�����U���[3�Ȫ�ɑ�����t�m>�l�kڬ�K�:��B!�Cx�\"*P��ڏ���pŏх������H��ʇ��(�~E/���6i�0��Iǜ���a�y;��==OwL���8�a\5����ʁ���������O�7�\6v�����⡋�����n�n�q	���(� ��B!��8�2yi�����;`g�s͙�T���S����1��k��{��=��3�.a����g��qL䘼s��fa��@�ɇ��Z|�%�[��}Z+QK��\�r z�̯��
᯼�jf���>+��:��p6�3��Ã��b)� � �-�Q0@��7G-�k���"X�@�0�L��hp�_�i�2�4�࿃�U�"[J%�"��(��TJq�)��Tq���UJ9ԩΤKiEJ#���+�*tʦҤ[N�5�5�miIM�M��R[II[)K��d΅d��*6��d��Rl���RE�T��6@��$�F��UD�!����<\EΩ6:��Ǔu�l��y�sͪt�Ѳi@�!Q�˧2)Q�AZ� [-�jwb���S�]�[S��'#������zs���ιYXm.tڭ�l�j�;��3�+����ㆧ���j�zqC��Q�f��C���^3�j���ʁ�@���K��x�hb��z��wci��;�ڏ�3��<|E�Њ�>N������dm��<L��P�\3R"9�*eqp�\��̈��t�f6_u��j6���jFѺ���V�^ޗ�ګ����1m���h��3������
�2��<�6�'������������������������������������
 ���g�o{�������`k�gZ ̀    h4���<��e(�  ��%DT�|�Å� DP
 � J@(
��I@�U$���
 ���EP( J�"�QA"�޶  �� �� ���΋��3�� /�	AE@
R���U]���۞FH i%��� � ;�`C��/�P��@SKFF�   
hW`�  ��/f\  ��  J�t7�`  �<�� @  E�YX  6��P((
�*PE	H(��H�A!!%���� !W�>�֪�    ;�#�'O�}�'���j�M�   U
U�ɠP@  @QJ$IQE�<�	��� � � 
  �R�A@��DT*C�o[��Ԓ���k5\XJ��+#$H4cY�U�
6E) ���ޔ��(P��G&���:��o�J7�k�1� �0o�U�
@X�@�T �x��A�P@�  ,6      j p w�p�Ѡ      � ��2i�FL #FI��&*y�dɦL�S�e1�Oi��2h�0�i��S�<i����� ��4#(�L��!4M3T���=@��mM�<�4m@  � �4����  C@  ��  ���"��d=�z�C#)���i�i��	�CL	�j`�F@=CC�`C	��C&&	�CLFF�`i�щ� I�D����A�1���(��bi��4� � �2#A� h4 M 4  �  �%(A'��MOT��44�<O�6��OS�'����O$�4 ���h�&������ML��S���d�=A�zF���z���6�@B��44�&&M24jm4z&4�h�1��A����&�L��� �O&��`L �6�$��0I�	�m)�ڈ;[���_Sbʹ5��}���'���B�j*�URH���5g׶`c�X�,h��&���@&����Pe�	 E��8�]���6I��Z1�nL��Dg�v�n%)qn܊-NoN�ec��q9�`$�[���c8��e8P�n��cV�0� �f�n8���(�4�.�ᵷ��'$(�`�8BX���H�$���+���:F�w^��kc�;��������d�2�`0`�ܦ�K;#e�w�W�� bCru���, A^)���Ùh4M@{,	W�OC�3�Q���W��}��]�h��F���ɾ�-��0�O"D���� ;�Z����~���2�іO�}�>й>����iM1��0��_8�/�������5�0,s	�5���f�kF���(�Qx�cn(o��6�h ����o��p%�#�|يڛbg��m�C������&��~g���i����A��K��g�3*����(��%��3��- r������	�Ft(l�"^�֟x���Q}\�Y���j�W�[��X���x:��>�}��I{ir���)=��9Noy=�~:��#�����Q&2�	�>���}�6�aӡ0yx2�7��׀�@	�TZ��9%+ C�����̛¯m���� ��{��<<��|,|�����E�}�RE]/ �����h������l��
 ؊�@a��cx�:��.�b��Qb�|^�8WX�xxs@�1�>���@ ��ʌ	�,=Ĺ�YO���b1ȇ�6���;�_� �'޾��m�պ�x���\�fǺw����"HC�KQ��:Q5��Pk��>�ގ�,������C}�f��f� �4��5�TNUFFQ 7���u�O���&5w;�|�nLeLw��  �< w�, ��٪F\H6��Lm"��5�L�H�;�$��A�8V�KF�6.x�&q��j�U�dS�ӡ�VʤDG�}@�7�ϟ���oԋ���fg_�BP�P	�x&X@2��8B�S��!"�-}fF �8�:la� 4a�O��G��/R�Y"�
���3��-#`�%�d�:u$��J��өϾ�U$�(�T�Q%<�2�f�M�P��ȁ8�~Ŏ�>���<��f��F2@d��"�&��w>�9(�����ٱ�6�/:�B2$2@p��jg����,��S�[o~7�XIǾ>d΃�z��e�J�4��)
�����E���c�J�]���!�S�����I7�Y�`hT4�$
]3iy��Z����p�M��0���̓c�2�,&n����>�`��J>�m�5+�.捴i���,3�B�F�-���R�^󣓞$|�E����v��UV3�9Pd�i��J�r�<U|�׏_�a�`IXL曭4l\#�lg�l�ٸ�ͥ̉b����߯kv<���������"ÉʲZ��&�-,� ��
���Ixr��C����B.�z�������a��*��ݗ�4v������e�y���3��9�tD�%�=ط,t�@� T����|o��v0At�����W.\�Ӗ��6'B DE��Q�ʙa
s86��%|
�~9y��HjX�`���XW
�	ƨۨ�e�9�Q�`P#M��+�d������������9��x�E���~�� � 9�P,�vJ,%!�S�x�λ�8 |��GH��z�bbb�,��9w1�N��xn<4����a��D�]{c�4" ��A; ��c�< \����s!�o>���4���>��3��k�za,`.�l�_��|��1�,��6a���P�����>��~|���t]�s�[}��y�Zg�!5�/"�nr��y2Y��}��&�@��@�u�����"�DA�&y&��L\���D�l��@���ࣴQjB�^N�BG�<��Q�X�R��ٻ����y��7p����@��#<�|��`S(w<cĀ�4�� �*�$! �#�����[�M9.�^ܼ�Rz.V�Kj=]pO�s�x{6����j#}�7N�`Ͽ��ƭ<��α'|ɘ�l��k�উL���=��,͡�~U���j���owq�ܴ1}���i�.:4]3�q�e�=��0e�v3���������Ƃ�Z���{a�-.�Y��J̎��$VD�RbUPȂ%��X�D� fDD �s�D�B\ؠ/'�8����]��[%c�o�w"�O%��DS�[��x��1I�N���H�w��4m˕d�&��V�3�7C�׷R ]���}qϚ�Rw
q<OD[]��,�%���Q���ڮ#�1��A�
f��ct���3p�F%�;öCg�A�n�Zwi�dFfh���YYU���=^��sc\�U�%p�O�ζ�.��#5��<!D��m��XRc5ɵ�=�kE�<7�Y��4J$Vs,��]&�ˑ8oݛ(pD��{�4�!��N.uMI9m���!�j։�}{C��>�y>+q�����t�mWg7��J�}��3�F�����4m͹�	sؗcV862i70Z�6�5��no�r�3��I�E{�uV���48�MI��<M^%	�\���D��!9r�jL��AL��"B��Gb�v�S��S<�j��޹���g��J�Z�N�F_2�����*�&��rc4����ΣV�1�ۡ�R-�|�úh+Uڃ0���i��C�{/>R�1����6�{��Ë�1j��:���a�C�����m��Q�׷hM�7�n5��G�W"�b�/M��(N�J�9��]������zut__M	��L�S�[�9v>t`�I�����D���|�n]v=����S��E"B]��^f��˚����Ui:�xj���t�y[��۬��k��I}zD���렽y�e��jG�v�u)���ٷ�^0�[���8���b�x���j��q��'�<y�-+��JY�3[�@���9��<!���d�ᛎ�w�ǎi�ܯRnͯ6!/ׄr�ms�u�9��O�կ]Q��������џ������<�6��q���׾����$3��O}~~U��pç~�˸�:m�<5A����`�Y#>�Y�wYv�-DK���"�}����������O�T
���/r۷���W�g�t�i��'�z���y��8���w<���S���d�Ҝ��s(~<�{�S�kG�H#`�,҂r ����?$��� �PU�vJ&@e��H��V]s�t�G�ȏ!;ڍ�ۈM�cs}��o��4�j$��t�D�{���J���%bZ�6��Yd|�lI"�辳�`��� Ǘ�h ǩ;:���d�Gt�5��X��a#x�3gu�/��Q����h2HI���0GtC�9��", !hH�s��5Ч3��6�l��Ӆ�m�ĬcI>�^�nzx�>J�BK�wmz�m:���+*wtҚ<�V��1P��S��<t�<k�����r�| 7�;H )Z 6���1���T\cx�:�^*'��t� �5}�=��S砋�0�Z��ک6�����������/,+c��zJ8�u�n+s�`�W�L�Q�m<�Y��9.KRe�(����ID���(��<��?s��J9t� >G1�^���NU4"=ށ+�9�gIvPcOg �:��:�Ӱ˺��#L7Gpt�d>W�͓,"�&�P�_��:��2d��0��P
H�	zK�.}:�ǌ�||�k�r�ɶK~��P��)Y�[3����1|Y�u�%~���=37^8s�v�y9���9{o��Ѫy�&Yq��ɜc�p��<���y��v�^��1��u�s6}lm���.ϴ��o�M��{��a�2�*�G$HP1&"���fc	!PP�a�.b�2
"� ��"�$��p�]I����� d~�I��M�h?"�k�p�.�s�u������u��.~o��p�]ZI��� � �1&���'���W�|`�<9  ����.u9������_����:�ؚL�E�3���Fa���?#T�v�:�D 車���l�_;����:s�hH+�p������y�����sF�#�vttvJ������O�!�ACK@��/���_���?����m�'`���0�z�1�ߟ���A�ݗvht�����l�q�jz�젊 �G�[��:9˸��uY����p�7�#��畓=�ٞ��Ď6�%�84`�=8W&�nD�]E�y��B�C�ap�C$O�+!vs�hÐ3���h���3�-V�ZOd°�/gN�c|7�W���/2�033��]ˍ3��B��Mx؋SÆ5[��n`Z�Q-��,��8����ό�J���ꓳ�؈�X����<(w���ё��DTml�����F�Ɋ�KE��0b���z9bml�kkrk����M^����{�!N��q9�\��v:\Kj�������\@��Q"�E�Ko��d��eb��4�5��ATET��I��\�F9��d���3��^�5�2#
d���S���1��<োO��}�_� ���G5rA��(���w�ł@l�-K�s������	��~n�s��<�f/��@��R$���K�I8�	|�?)R�ت��J�~R��p,Ap֢��j�%!.��{=�s�[��$X�;Q�Lf푪�~����xPVW��)��x�/9:��l�[e��S�6�j<�ڶW�㢈��o��δ���T�5ƻس��盥�7{5�tRMg�7��
8��qOHG]h�%�Jy�.&��8�GX��+P+4m�B�Ů{�n�j
�|�ǜC��3*-��۔5�MB&h��P:�H�-u�9ͧ����N�������R��" b	Uba��K�9���=/����"4�A�b��J��M�d$���R�ʬ���Z4�[��;��.�B'X.�������n�42�[aPiF��n�9%�[UV��K*�P��A�b��:D�XO�|��.�]�&GY哻�&;8Cm?&^ѱ�ֶ�Z!���v���:��ړ�J��zš��`��Pi��v*���5PԒ����{��_I�&D_.3������!�!�~N��Rvw�y�<}��sC۬iצ�^b�(OTE�}�'�P��+l�*~0�L���7�/�\���2Q��ݼ��C>��:���/	F5R�r��,��C�3�}��<�E+�\�� ▄���v��K��#0pP�+(ȩ<b�DAAO8���"ն�[�^�8�(H@����Ӛ�j�{l�9NU�Ǔ��w�������<M�����3CkAH�HQKJD�0�1�4��!C0��R4�Y�t�|�ՠ

�K5���f��4�����f[+k�f��X��)���f((�"��	��V���A��y}�����������g�#ɢ-Cj�6���CSm���vvX�.�϶�ƥ��Զ�iN������J��*V*ZY$��SJ0dIiaL�!(@��� ]��0�t��O���6z|��i�P"�IALA+�������k������`�yy�s���n���*+���"$S����n�oWe����Mjh55[F�!T m��?�]0(0�T��9\	��j2MV����j4��]|��ZKL�4��/]��F1� `  Ǉɏ�ӛ����7�{�-[}\im�w����y>|�!��ֵx|���m�f�lq6���Q��8KYjn62���=����AB�(�ڱ����~g_��v�����%�����+��_���M�؊]}�c���[��D�=u��鉃���~F�7,a������;�_�ڬ�_��%�i���|��~�=�C�͏Ӭ�_��g�A�g!W�����_����'��˞����'����uw����|�n�I��t��>�+�<s��t�e��=��ᏲX�6�Aa�/4�%>���]vGf/]��<�^�������H�l}�K�n����:}O��/m�/b�<���y���YW��7D����ps��'f���ɫ�����n�7����c̕r�ZG���B��㾏��#� ����7;�|Fe���T9S�Anϟ}�ޏ���fwLI��]��=�=/7ε���2�]���	�9ǔ�|����������-_j�E����g3�����%�~E>ﳯ���R��ٗ���Z{��Ҭ�{��N��C���MޫU��~�����3��|�[���������Bq�F���|���t���m�_��I�f�+�ð)w��P]����LϦ���O����$��U���
�,�L3�c� ��D ~���7�X���W�_�UI��J�@2$��!�"���Wnm��-��d��%2��{�M�Ʈ1��l��{����Mϡ�9�ѝU���a�ѱ���O��e������;��[�� �M�8=Ϩ�Z��v���de����l*���鴸mC�_j���4�@�!��.�FK��8 `R���D< <�0�>/�������9�?!��Z��'�dcՓ� ��Aِ�s�`�1�w�(���01���!��i�������|���c�?g��ڴ�ֿ��o��&@��z�K��6\^�Hͳ�ѻ�loB3�� u)�y.���%���6qa�q]�ϩD������� A �˰q,�������{� ������>�0���_> �c��ޓ�N��-�z�FR�A3i�
ax� (H6ʚIH  �03���!�(I'8�%I���(m9 �$�6��y|�t	8�_�oJ�@ |�L�o!^�6�	XhB�Q$��P��Dk�2�FA.�
/�s�ο�ԋ�� �?PD���1^�7�[��98o���M�VW�iԆ$zf�@A ��@I5HC�V��gu� @
?����HF�\$XB�@ �  � �M�Iw��t�A�O�rQ5����\42��p$\�L+S�����yT�2��^Ι�xƉ/:�� �P<�  ���F��#k��.�Wq��5�h��$�f��0d�N^9^   x@A  0!߇�n���j��ࡌ�C�g���99d"�3��]�� �M��oM�K<�z�*3�LQ{��� a�9?�/���\��D X�^1󣞕�D���I�O����c}����	2S��<�&1���HLN�̸ۼ�`B�Axd$A� B"P � ��@^޲!��E�9�f�Ef+� N� �;�ŢRD�yd��� �H �������\u��FA q6�${j��,u��1�oCw]"KS�щ`%��������"�dGR��l����hɭD��P� �)4*¸zǷ����D�DU�xHO��<���z��~���`��?S�}�n-M8��>�8p2L��i�x�QJ��bŢD5Y����Ɖ�Ԛ�Ti����e����D� @�HF�j����7Et8@�¡K���~��c�#s�]U���9�����M��>�+��G���0k��弾�$c|Z�$~��lRIօ����m�+�*�, �/�+�a��U���R���A F@ � ���n2Zd0D���_*R�E���3��_`
� D � ���~"�R��q��n
m �G�8����ΐ��L:�6��`�s�$#E*��s�0z�O'����}�72���N<�pf��t �    E�t`  GXd���ɜ$�1�	`��5��U�[>(7et �0�[͚pA  	S�0��\w����c����Z����;��l�:��ƃa�Ɖ�t��N ��  f�gB 4W4c�N�-{��O��7��~��٪��c01���1��t�#ï��M��S/�b�,y���H�NUF@����F�"�`�e]�98���d+t�)�W�l�<���h��P,�䔂�    7*��,ȨS AG{���J$��8���Ӧ�����<}�&}�2KN�� ��"  � $�:-I��뺤�:@w�&tz����{��꿟�� -�`���&b �"9I0]<aʜ# Bw ���¸"B)jê�c���个	�(�S8��C�1�Op����3���`@A 9���	|��@� +!d�j%5���ű{�)��!F",�M�aRi� �O�(%j�bC\��QЬ^,O�) J��Sb$�%���Sc(.ni�����%&��$�	��w�@�$��/��$(��H�u�RAA�%~���ޓd GE���������%:k٭�[�u��w��� �I  ��DA �B�I$z��0�	:�R���X#h�Z%�a5�t
��D�  
�JJ���5� �  �Ba�=�e@�&S-��"k��Vd�@�?x3�mg=�׵�Y�(�&E,[�X� x� ���``zy�������'���Blޗ�١��k��s��x~L$��M�7  ��$E�4H��%Z�u�?�έ��ㅕo�,�>�]���`��O�>�`b>�_�|שEч�`   ��56N��X0�*���y�4��̝_�@��  ��L� |���� �*N�"A�Ʃ�Y]���PG�����_mpEMȘ`e�) � H}E��~�J9�Ic �8h��.��uo�32Xቾ�ڭ��-�e.����v�:A��%�Ĕ��2�/�:�,��@[fh�{�E�$�ދ����T�A A�x�^a�	d�6cl�x��S�3sk�-Tt��Ia�Ε$�$#0`>~ƍ2jPm\ɀ '��� �Ǹ� �ΨIrD����/�!�窡*�y΁�YAY$���	o�P�3�%d�Ct˧]C���k$� A[h.A7�U6����i�Ĩ6�1�G��"�f�T � ����s�� A A$�.���(��>��8�-����e��,Ti�|oN^�4 �v2C$S�z�I��?o\�nZ'���4u�{�o�~AW��ϷOq~y�W}�m��'�Oue��O���>��c����B"%�`IU8�%�	�y��z�F���ʼ w.X��H  <�`c��q�M4a�v#�����oR���ϯ����O���{���^�Fo���9�X� iS�5�|\�/1� �R�$^���`'�yʼX�i�y�XW7�MTv��^��� u��D`A ���t��i@�;�&�*��+�R�� �Ba*��g�# �6���K9�O �t2��&tU�֐i�DS�r�Ȱ[��pu^��})��8�S�K�F���,ɶ�1�xP�a �` AX '7v�G�����DVX�q��ݩh\}�0\~QA AyB��wʀ� �3b�W@&�N/���
�0U��_�8��bcNz���� �*9-�4��f+�)�{
'���8u��N�*��!   ��%|�%P���u�B��k��C�:� ����9���Gbb�~�u�S�H4�:Ì(�]9��:��Oe/�dD�;q�*���M��tp�  8٢�Ru�	�O?���\L$��bNyz^��d���ㄋ���I%�  �X�-�M  �cʓ��&輲)�Fs�9rSfi#K@J��G�m��Hfa" ���"��P�6� �ɻ�@�T�I�I�{�<h�HW���-"D����;L��%���t��@A B�y-Z���kQ '�ir�t$�ȇW����1�0�l2^��S5 ����L^��
@k)��  ��H��}�zi]��;m�� 1���w�d� �o�`c��%2�� Bl�Ѽ���6���r`�Ȟ�  A @ @Y��l�q��Oy�ћ�Ϛ.Íe?ϙD5�DT�Q	��!��r���/�y��Ǘ�wt��Mb��9�.fa�wn5P�-�e�k<:˛��Қ���ڽڳ:f`�+-���0۩����yƵ�jY�T��m��0@��ޝ��sF�8uF�������:k����T��ry������љ-W�S!!k��Z#H�[�x�Y�\.�t͹۪&��զnc�s[�bS���Ś��ҍq�kD�h�Xn�ۉ���fs�� e�Z3H%��n@�$�Aii���	!���-�&��-��0 �1�U�Թ�t�Nkk��x�֌�wm�lE\�)16곌�x���M"(��U��@��U��Ɯ��
�ShPk�r�I��M2�'Y���n6�q�#��Fj�z��7B�m�i���ŕj�x��UY[w8�p�Y��e�fr�s42cD�fm���KW�
�����$�u��1, B	&�ԧK�F���ۭ��C܆*��حR�)S�p�z�qh��Kl�0�BᘫR�r��i�̵��sh�z&*k�2�73%5�ju���E8��8+A$�e�&�0�D����mi�n�r��5\\E��`�"�$v �%�HI$k��l�My��&�`����NP�w��`-��n�f(�E!5J�8���j�QHԘQ���&�	#����JQps-�rsn5-�[m1+�k�.V��*�.kI�VIZk)jӨ�i��N���l��ت�cA��	*=#Dvڗ�k[hu��d�̭eq�0y�������w;�D82�1=�R� )h�B&��(��,�jD�[%Қ��5����f�1
#L«�k�*8ƈ#����d��!��e���B6��W�r�pLX��n��2�g34��B�8ʊ��ݷ8���eJ��Wqy��5��Y�׏Dq�e�ŧ3wfP�)K҆cRR���BI"���l�A��X8�-l��@�Pt��D�9P���i$Hƃ�B�`h4�.�-�wnN6e|$��諐9��7HL9�y���vNR��G$��O�ݕ)���6V�$�� 
@ �$����wV
Rio�UxˌF����L��d�PIV�$�.�&�-�0μ}��-�[��q�\�rŴ.��������ԫw2�G����\7.���e[-r���U.N�\�;e�Q�:�e��u7R�j�[�ڼ��Cn�2��F�S�iKf8eX��m���1��˃�I�LDs������*�����Q�(�֣i��v�V@�B,�ME0�,5�Ɓf0Tk��%
�̢�M�ek2Ԫ�^4�-(ښ�F\���TM����VL���c�;��Ö���V�0���D-���\�U-�-[X��zaqEKJW�¯KlR�ܮ���G3�5�tQ�Ն�T���C�����m�i��t�
�X��q�,u���^Z�)Z��[X8A"��A�Y��$T��53��sz�M�H@@��b�L+&���!�Mi�F�eZ���R)u�̒4�!� �[��kb&3X�U($*��Q˜15��2���pˎ-j�c��냉TKJr���Sm/r�����6��++ĜN c��CFR�2��Y�\������8IdV�2�	�y�-9���ظZ��u�ne�4:��+��x�˵���ݤ��ѡ\�^7Ȗ�՘�L����%t������%B�d6%�-�ف���hb[Mu�YYG��bM�6Hd��`XCH8��X�M��(���p�n�܊&:��f'4����ŏP�]q�������8��c�f˖�,����"%ax9�q�U��Vf7�E�9��p܌�i�Z��m�#�a�pqp����qe�b��ݳ�\G3.�X�u8�l"����j�`2�%�NQM�Q��J�������R�;�<�1�)�+5�kSr�4������h��)kZU+�W-�/x��1(�*��QE4��DPU㦧c�!�ȴ���+�^Xq�N[�˕�Z�Zs.p�0\�Wu3-2����c��6Ŕ��TZ�h\��Z��b^��Z��e�̭(Ws�P��-�*��e��a�lS2��,�ˌ�L��3�t`�yh�Jŧ-�4W�LR�b�K�*�����9�x�i�\Z�����R�Z�̻y�\��k���^Y�����KEe�2�')X���na����-b
,�*C��q���Z��S\�K/Xk6%R�0�*e��1B�*	��[�)��4L
ʵ*�j@�H4�ȷ+�JӐ�-�[]nM��5�֤�\h�yi�5�����9�m�ǘ6�u1--�Ҵ�c�y�f�A�7031�����"��"��i�
��B&I�*g�0luI�Q�'0�*e�k�cF9J"�ט\�(kJI0�h�Xh��k�sp1/n<��V�j#U10q���z�&h����c�h�m*k2�N4�[����Vsi�v��j�ѣU
�YR��ǖ�[�X�[�*�q曕q��q�ay�U�]LakW2�\�-ܦEm��(���9f�7pj��i�F	+E �b�l��,2
��4�!�l��K"��,M�%V6	0�����i�eBʍ��۹E�g32�-b"⅒$kN��D���+e�$qƺ×�7&�s����ȌEDmY�)���ss.�J�is(c*9qy��]�ԸŪ#�-5+R�sh�ا2�)S]I�c�o�q1�ƺ���\N%E�˳�
ŪǗu��ܸ��-n3���֡P�����Q0rS2�r����9Mң�ʢ�yLۮ��*��'L˩�0]�[]���[ĳ�Ŷ�q��n�X�XÍ�qC� `�4i�LL�R+˱�r�/�-�����%-]smM��[mL��m�©kI��2�ݦ6�����u�)WR�W\����.�r5m1)mn.�1�dl[Jbm��&�Q���&��5Y�6�,-���DEt��҈�B��h���W9G)8�`=�#bc����Y�5���{�మ�e�
��R���e7"1 �*��m)Yw�ո�;$�(�� ~E�&,&ձlLbS5J4�mX5P ��ݷ��>�n��H���'���{/���̟�7�����?��{�� �� @�
�yT��?��;N����4p�6�c���/�}�m���vLa߲��=ǘy׮��0������u�@  ���%��P���*��I!����e�)hj�hhh�(	")��

h�����������b���X�`(�H�)������""�$��"���*���!�*P�*�"J���b��h�BD>�6[���?���!�z/s![]~���X[V>!z���%��Am�ˀ�Ś~�r,8� s�&{�	C��j���&��O+#�<S+s�k�~�!I�����k�5W�d�MaJr��|���5�T�zO�+s�T+�|}hD.
fPs^�^<ƿ͚v	�!!x��*�z���,\M|�����Q�m�i4��H�|me��oq�Q5[b�zZ�˯c,� քc'�s g�&�'h�6Wδ�/B�e�g�ӛ$�t�-Jf[
Ɵ2HK�MF�٢'�K8�c;����a}9Y,��F|�Er\X)#�n����-7*���re��̼Y �jÜX.�|�쎴�:*�aFV��O5&P�֊R=-۴�����,Pb��͊P������M�*jmNږi�}a��0�mKTQ�O*�����¿%�5��\��r���I�uLyv��L� ��9|k&�9�Wc/:��c0�T�~�2��@X�wp�6�dF��A��n-L{ۏjv,Y���:�(������Ӫ5
�L5���,L��˻ev`����fcm����G��(_�
�ĺ@�� �F�
�˵c�b��`J΢���s��L�ɠQde12����l�If����9�I|�D 
����{��U�@ K��3�� ��
�:��-MVj#� �%�ӎB~G��WҨ���C �D^�o.p����z����v�=�˛����v���:/�����M�����������##9E;C7����j%���j���X��ԿW��	,�y���R�UȊw���T�6u~$X�+Q������?����H4S��Y����M�#���$lʤ�/��	�B������^ѓa�R�wt�]칓>MvǇ�<��/�O	�ὬM2v=ٯ,��YZ��D�0vԷ,�6�K�%uC���K�y4�cQV^ӥ��\���>�BE<x��w:�R����)�GNsny3��=�Ի��"�9�,���Q���gNR��Ĥ�]H�e��\:MM�5/c��n�ea'�qTB��b5�ߐm�aT�:��_!��H���n��`,�JD�ެi����/$���E�m�O=��=�(��<^�~E����T���3[/��[����F���\��u6���1�T���SrbQ)<�'El�s�_�M#�WE�i�o���:�Rs��!������DG���_-\I��cw f�U^n7}�&j*�p�=�y�+N,����*�w�� �|&>ᑹyQ��$�m�&)i_C�Y�MG�?�wc4-��c�}�)�LR��u��f�`�|����@ԥ�1j���
��8�1�H�v��{0�<�uMT̙���wA�
���]N7�F��.%~%�1eGS6e@5X�p��˞N̫_�.pP�q.y�3x�2R6Mpz���[g_Z\k����q�EC���<�ttK;K�6/&�oz}54����ɡE J���nA�gȹ��}�o���[�c���Ѿv���ϧ�om?W���D��sԵ���	yB�&�bΣx�Zݩ~W����3��u�bоaȞ,)@Z�xcO��m��x�n'=��<?��<_	��&2�(X���_�w�!t�&�b>x�����_�6W.`
V*ȍ�[e�c"֙��&5�-r��pƸ)[hej��f�L��D0������c-�ĸV�s��1$�"����,�fJ.V�[j���E�Re)�Q(±s3L�Ź�,P�69�8��LJ� ��a��q��U1�ƹ�[�T�-b�\r�Ĵ�qs�-�qZ��E��G1���D���)��B�^n�X�ٛ*�Ls ��[J��5�W��扲^G"q[�a4ӵ�On1�
%vP�G(M���̨������%�!�)�*��dU�!>���
Tyr���\s�3�ՉE����̣jV��j҃.e�婕e��q3�G.8ܹJ\�\���3
-[V�3��p�\Er�.e�e.c�m��⸍�[����5r�j��#��.&33L��щk��c�c�31�3̦1�m�`�.e��UX�Q�mn��"����!!m���H*��_G���S��N����E.�t��XT��d�)���!ۤw�ToX�N���ߛ�n�R� �Q��YN���zo��z���.ewj(��#�U�f:tPڐ�}�.���eu�����-W0�w�:��L[y��{�Y�!^����Dw��]�wi)�=��鋾�u���)j=�w�{̉z/"=�_8��Ocxo.����
>���¹NGv�y5<t�zT�S�J��N�Ox�fV��XZUS,��R����(A>��3�:�����b�,^y
/5���.�^�.��Tz���׍W�{xQ�ry`S�9@�U6{L��&���l��<���a�5�q�ޏ��F���.�P�%]�����.�޸="}'Q]^zW�EzH���������_ h�ʞ�S҃�H�zӢ+΂���y��U��%����P��ޓv��׷:ӽ��s�z�7qR��^M�c	� Lq���ͲHB�HeS-
kK�T�(B�,�d	�,
ɻ�ۉHy�9ӯC��q�!�]0��®!OQH��@2�������������8�3��>�2���ۭ�v�3�z��8�������c��z����f�����C�T`�91�O�����@ބ�IM��,�	T����~����>G��3j/+��h�g��������a��wG�̀�1�s|�<�&|�;d>�G���a�-$O�}\ #�,�s��4���3�����������v�.�s���ƻ��,��< Ae�I���q4H HIO������$1>�,8v {=K��W��L��������  �R��$y4�Q "��?�����>��������q����+>�o������Ұ�%�A������7$Ma�_������4ڪ�Ә?3�A�Pu˶s����:yzB\���W5IC��� ��RSm�;/��T����ǹ�������B��u��]3��^����������f��.'�@��"ZuViA=ʟ����_�l�Pos�L�O�d\!�ɗ��A���4J���sJM��2u��e�{X|�;t�����?�t���~�jT�����mR���ɹ[L4�œ�g$�[`թ�%W$�AX�I*i�+S-�+,6������b�V6��"ɝt�]0��DQ��4��TU-T�UC(D�E$D�ĭH�RД-%REQHU(�2�\J�6�m1UlCi6*��mD�b��#iIH�8�DSiSjW�!���y��"�&����߷��
lN!�S,�e����J
�Hڪl��M��6T�F��m+bm�+� �U�CiFʫb�Tv�qX�_�Jzn�9!��;��7g^�'�Sal-�b���;�#��d%�T�e+iA�	9���;�t�9�:�u�G]�W~�����A۷]�MR�~�%;��*�m퍀ڨ[l�9��̤�9����v�bw�m*�m	[$����5jA�Tt���tU�s&�2SdW5T�Hۦ�Y��BT@�6�aXp��n�&p���TF
-�Z:Z�I��pi�v�7�s/�RԸm%���r-r��奪���x�m[����I��
#�X�̼=�zӍ��ܧR�L�j��h��-)����k1;�#�9LE6�2���T��`�v�ヂ��Q�b�-��]H�Bt��%(ㅂ)Dń��@if
^�d�ޥ�VH �{�J�fT.4E1.QWYK% ��Ri6���tL ůH�a,�`����
I)��ԉh��I$f����#PF��ajh"�'$"��5X*�,0B&���P�5Tp�KM��$g-"*8�j�ZT���<�]eM�m%���&�{�I�AV�	+Bu)� b���q0��0�8��ATH2�e��	�F���Ng\�VѶ�7�f9�B��[-[��F0�8��	4k;�/5-�)���M�S[��g�f)n8.�E5��[�nh=��f�*\�^���V
aː֢1u3.�ܮ9[���Y\���r�kT{��l�x�I���g�S��=�L�W��Z��m.*%�˹s*Tj�Z���͗��e���S3)k�W-[��#�h�8���!��k�s1pA����w7r�fSj�,ƂAS�[hhD�(X6k i,ֲ������Q��*̸`U^��x�TLq�y�b7e�J��0�@&�����Q�"`M��f&	m��nk���an�э�9��/t�J�ܩ�a�a�N,h�,�!ȫlF�$����^%��8*���P���5;E1��0s��-��WK�yxaj[��*(ձ9�d0T��-�;��YZ���q����ͥ�Lq+i�\E��F��r�"A�a!�Ј��a�.Y���Fԣw;p�jZ�E�����r��w��+��+���4��*Q�D�35�56ّ0ܮG��p��܊�EGZ�ۧo1*�7�:�;�Ì��ۤțWpƮ)�uf�Է�e��2�L۱ik{������ӭ�\ͺ�"ؓI8�5q�D2!P��Xf@��p��p'5ƛ�j�Ie�����J�����X��0��3
���qJ7��H�IP�J��~K���S��C�I݀��b�IyIX���!����~m�;�W~K��P���@��x���c4Wl��w��듮���@�Cj���&� u��<��<�!�������dC��?_�<,�5�*H���uԿ�F��9>ÿ'�`��ᖸ
;1Q�G���E%Ms:BBBb�1�"�v�m��b؛202�iF��b�b���� �I�eA)Q"���B���b��`��hbrPȰ ����v�2�<m�����`�hA�
�����L�����'�^O���I��B�������I'�k�D��j�;����Z��ߖ��׿��'O>���9x������C����f�?��u�C����������u�g��=�����}H�����t�o�������3�@�I�nze�'�[��o�7���}���f*ȓ��\�d����,���d1#,J�醮|NN<9����˦oCa��ߑ�ݾ><��/�0�4d_ŦaS�ٺz���=}QM�E6".j�J�4(�j�ps��Y���X���J�*F
R���
����-�H9��ڤ���B�UmA�I�l��RM����	6(��C'yV>ֱ��+�YF1r�!�w�b,Kcj�W��J1a�ܷZ�C���t��98U�L�OG.B��
�S�n+�	���7,2�Ap\�8�J+2%Ads0�
��r3�ձ��LeQDB� a��(�Xj��U��m%*��U0�V*�U����Z���1��:Hh�C�	��V@Q	'I�1�bb!�
���[eEQDV#�A��(�U����J�R� m�E�X��c#��@��U�Ld�6�h��U֬L)MJ���1��3a�Rд�*i�(�@���6I��T+**�b#mb���U���Ab�SDf�*���������>Gm�����<~�����]&�gU�u������{8.��x?���p��C8d&�����J���KeQ����`�E,TkTc����`�9D��|W'�o��~���n|�<m�{�yK���|��UѝO�1Q���c��vX���� �ܚ�w;�_�C��{MU v	1�1'"�"d�AD"2rإ�Mi�UQLj�1�R��
�Z*ʅ��0�Cݒu�9��(��U�
"�)`�Z(�* ���Uf�b�8 �k��i�~s��_��eo�t���+p3�*ڭ����?�������S,\��M�&9���[�=��j�ۧ-\���T��6],2��^�ͨ�Q�GtC��:��àH�~W�R�M���1.qE�2/�և@��fwu��E�=��:�XFjɥ�Z�l\�7��Tm<q���
'���C~)˿�$0_�-2�Wi얎�#fז�sf��ڥ:ůu���ް0��N19p3�l�k�h����.�*7�@I:l�I��.16sҪ�6pi�m�'"��eŢa#�?|ֆ�BlЧ2�aX_�ɋ[��
kּOC�h��X�>��"�%�x𹈴�h\�D�[ >aݹr�q�٨����+x\�чd�[ˡX��t��==x�7�,��É����*�1\���X�F�*�{�^g�*c�V寛�\�*9��:��C2�Z��h񼳨��9\3.}���cЙ�h��6SB���E�;�On�1?L��3B(o�tv�ņ�c³��-�o���ѻ2���Β�jF�Ѷ�Ya��[�ܻ��يU%i#��p�*j�MGST�V!Y�j�m����N=|�IՇ;�$�>lc&k.\]DVL���.exs��r�n�Y�#��km���%Yv
����ɩ��^V_j;vӺ]U���-���_I����6-�M��BV�f�q6OʶMj��K�8��\VC��b��d�2li�n�ja�B������=�i���Z����43�����ց��0����6"�ɱ$�8��9��=�v�w��������`�[�͆��2����}ԢrjT�U"��X�F*-�Ab�IUH��PR�Y���q�N���'6���C)J����,UDU\Lf"(�����+��]����bd�H���u�Н�z��7w$�.8e��eb(�EX*�DƊA�qj�;`�,��N�'d�Abl�Q�AU��"�*���"�YUDL�Z���@��#	]	ᡪ�"�ǉb��+m���1��(ۙ+�,J�8�b�1�J�P�8q��8�"���E*J�bT�e*\�;>2Ϳ˚�sp<�'������w������x��,����������4����	�X4���mEQA���\�4SK΂ĸo�|� 0�S?���mÒ*v�g������qD2��/�9���&͕$�r��|�IۆE]O�B�A��\䚃��+��9L�T���s���c�E��Ԑ@��
?��?����w*v4Q��D�OהXX}��]�
�	4�&��['(;��T:�f<l?
��i�)�d�-��� 8�v�.���Nǲ�,��E�m.�2A=��茊Q@��"t1mІR�0��l�-H�Cȃ+"x���h�4&$�7,�j�75ک�6�n��.��᧨��c���&���e�6����m��b54G`/D ���!�<`�XВ�+,�܌)d.�K>�of�HM�`��h�e�M͔���^�5�]���Bl�M�3�K��,n�c ǥ}�&� #�<21F�n�A�dJ��w�ʴj%2E���R�Uc-��5SfZ���]�՘m��������b=��׌wKV�!Y�;�5����KCH	I@�H����@��qQQQq6(���A�شH��hO���d�@� bB�LD,b��R�C�gm�I����X,X�uE��(�MDI�TU�6�EX���`����C��
��ԐRK��:��F""����TbȨ�*�H��Y$��0��'�jT\`���S���Ix�;i��R�J5(��Ak��I�%�d@��$�vجXVT����d5Nw�(�U���I@�)"144UR�H4���PPT@QH{5`x�aR�y��-��J,�����1j�C�ɔ&$;��=*X��Z4��J�,%�X�֏�)�fa6[V͊[�[l�[N:���Q�k��XF�E�IE���,s�.h3�NsC1��"P��J����b)
�pL��T���r�eb�XEJ�2���dF-IPXTP��B�iث �KR����J��+
�J�2
�D*�-jK�(B��kbZ�-*����-Z,��B��a=���?���F���3'��z�o�����i�3-�܅a����װ�H����~(�������Ҷ!Y�7�[/���<�>��_� G�o��5�k�[�'�b���֞-�=#����֕��p�R�4��)6�3a@b#f�YY$�	J�eh�JŔ��[J6�J��6}�	��"�3%���I�&��Y��)�TI:[ Y�]h�E#6��H(u�b�eK��
���9�(Jj�J�("J$Ě��2k(�X���):�k	�
���*�R(EaZQ���
((�1b�hI�����CP:�2)&�$���#B���&���岈�����5+Xf��
�U��I�nL�ST�@P�I�=$�ݳYX,R
)R�Pb�Y%BI%I$�0�u��֣"�XX(,�Z�����1$�NP�$m�#or���A@U�`)���RHAp��yh�"�$
���0+1
�k�8�ȈEZ�dQd!�I8�	2N<--�AT�����,	PY�) 1�;`a�5�$�%H��F(J1E���1Ɯ�sR:��]�����:�QaU13)V*"E�	P&��
Ad��1�a1�֢�J���,�! �&&"�q��Q(((G-T����HId�N32�AaX��"Q�aPs�t)iTA�	XHT��!�$
��	2��d�+"ZAV**N��
�
���UQ�X,+&$%IIRq$��q	��PPQC*������UF-�QdET��ے몹�t�l���9�,"���du��(�Z��E������	P���H)$`a�RLjJ����X��.5fR�+Z�X�� �$��e)1���d��2c�Z�"�EX�3(���UF"���h�N���%ݪ蚶M	�ơ1��1$Y�Am�[h�b��*��c��M%9�	)M-�U �Ɉ�R�I�1
� e�\��,���V(�R�Qb��l�`�8���/���9�Lw�Q�+i���K����cFi��� 
�(�$ʦ� 5TE�I�E
8E���g⒨X"��f��[d*)m�"����cl�eE�"E�T.0@������}������漗9�����u_C���Ͽ��k�����.o���C��[K��^��E_]��Gp������O�=�Y��e�Yev��a%A>� �2Y�'NF4kSy C	�K�u>_�����<�h�Yu?������ٶ}_-����o���t��l_Wc�6�[
�ڽ˟���g������W��5���*3T�4�<���a)�$���C�M>��\ %E+(��
�{���~q��͟��3�N���4��r�S���/ۊ�����C/���}7�1_ͨ+}�y�N%��8����H~t������e8Z��o�X{2d���(�A}kk�"7���&Vدz�'MI���Č/�}:�ےW�sa�u�߆�uw�wg�E����jC<�\�A]T�;U��;�Qm��̆7d踱��)+��SzT̓e��X1��,T�m9��$�ٙ�Z������2�3���w�L�VXZ�cc�퍜O.s��_��w\Xj�	F�$�[�i.�pl֪�,X�������gx���8��I�f?�H�{�ۨgm�/I�Ku��b]�n�е���=�r�&
�$dzԐ�
��z�̔�gv'Ңx4i+*�Ő�qmY��k%�������)T�h�Ԑ��mX*R��nz~V��̴��S�� ���po���6N�Z���c�����q~8�Ӫ��y׿� �ǖlp��������[vhߣ�J�nڤ�21//(��.JWr8P���^��Ֆ���W2W!��������S{z�hd�x��Ʒ�RK`-��F�89���oB�x���}�,�4��a�`��	g�"�e:k�T�vB�~<�t�jtKͭ�6���p����k�$ُ�N�!ȫ�͵2���fV�N	n���qɽ�N�M�p
4�	*rs�V�u�����oG�lQT"�z�8b�8
+�A� A�w���O�����tyNx[Pj;ޚ�FJI-0e�e�0hƔ[�PN`n�� čH����8�/�Tu�Vu=�޸�ҌD���?����T�����Ī	�{ښ8�qg��� ;�,�����`��J#��|�*�뒙�	QQM"����xM6߸�S��t!���D��ʽ��3����2�9�WI�p0w�}QC\~���FL6�Y��מ�3�}�v�Ɂ��V4ޣ)����A�����H����VU*J,ؐQJT�1�|�ܽ��o[���O�`�A����'�,s�|1�k�/f+\������pi˝2�-=T�Z�SN�0�K�av-�5Dl!^��|�-Z	5Nb]i�.z���.�踳O�� �5�,��p�kr�a�yi	��*7��)Fi�K&�?R�!�)}�K]v�A����22T� �}�Ώ�{ѵm��_V�e1�3�S�JƗ�Y��E�v!�ԧ8�2�~�8����.ؖ^q�N���N;��m�)�� #�FLD x� ��JZ��*��� Z
A����)))h������""Xb��4�S��zp{Y��_��Y{/���g��>���w���1��.���H�7;e��Ɩ������j��sk�����h�?��O�A2maW'`�Q.h���ϖ���������a_@����hߢ��d��l;����]�ʨ��<����%���F9��7�e~z�5#�alfĭ44���A@RJ�A$�Q�R74a+�P��@y�I����(�� 
i)
JT�sV˝YۣsSMj���-ʝ'h����������z����>[�{O/�}�nk�q�>��<���'���_�^��;��j�� �,����m��ٗ&�e�Yhf��ٰ�Ж�V�m6�6�lQ9��4Tڑ����h�ضD��W�ʕв��r4b�H�B����c�e�_5�?��v.�����x���s��zE�w��[�%��W�;����*��(1�YA����=���ޘp?{�{�{?e�q;�wfs+���>�s��k�'yg2�J8��:z#��H �H Cgܑ�[��{�����=�(�t���kIw4e�J�pa��/C���.��Kz?D��J�c��W}T����{]�N�������.�`mi����ƊK���5�ݨi����0�[�MJ�.����=�'����ݥP��!���/=�������+�Y�rP˲�m����c�Xw���t<���D�H�;}��d�sv���/��m�_�S��~	.X���d�����ЉB�$��oq�~����K�m~�r!��y���'$[�t3�Jíïe��%)ft�`���������{���������/V(7�wf*_d��V�[�eBz�CF���ӣUC
Uޥ(��
�ғr��qSR0'�p�5�$�;��igG#�.�1�S8�Uӕ�����\��!�a��;�M�?X]��
E�,������g�ceҕOj��E�+M
EW�`���́�3$�	�:��g�t���o��T�Vwa���#�Ͳj��Q�	�dc>��I�v75g���rp��E�e5v��D$ӟJ��B�ʩ��5 N<
��)�4�J���Q�5�
M6��7i�سK���nߕL�����ԥТ�����k�6�z���d�˼�y-��<���.�N��9��68�s�]��s-͹v�����o2��-t�H��\�&�g��3a�����I�
Zõ>X����vRz����c4���������ո����lpRe�)Gf~/p�y��ͳ�z�E�T��5_���כNr`��N�ظ^,r�h<�
迶r<ñsd׿M�6��{��)�4l�>6����h�R�  �fB���\''��9�c�ױ�e��>]_S�])�p;�I�wiMF���w����t�@}�S��W,�I���r.}T�_�����o܂̉�_���Vi�	~�hL�o��I,Ba���1}qt��7�d�#�k��	���j9hEo�{ojߟDBt^������	ݬ��c�c�۩W9am(.��8�Pz"X�OoyԐ`)�	���zN/bΚJ��J�F\�|2ݼH_��Kr5q֘tEY�V	�k��h�'	`#2��h��
�W�<�"�0��Gx�Pl��G�j�R�q�$�D���$��	��M8"P�V�o	�	!�V	YY"���l�X����h-2v�hkL
�����Bܘ�d1�q\��34aP�Հ��qƲ�q�ō�=揅�c�A@�L40�*sMH
=t@�Ŕb��ʉ�A���xm����{�n	�nEe����#���'�
� {ͦ��\�9������ ���RMp>zt���up� m#55%#�KS�V��q#��&����^Ö	M$SR$T��s#�sa��kZɵ��!H�"�`�d�,bDQ��
� z��w�_�y�;�m�?1��>Ǟ�����ǟ�����O�wn���^������?V������׻�����X*�g���؅��l��!��#�Z��ʲ��d���HHQNO���i�s�t�?�xñ��)����q�O�n�n�O����P A 	 ����Լ���cY�>��U�E�x����py�*�}-N�Y�T���ư.���;����	�����k��r` D   D@�� �+��l��V�^!!�y���xt�w�����ݹ{&�{�R�-��poeVR�1X�!�C�U���}CS��wM"˫���=��Lv�r��7���͢E/4mW�p���i;�}K7�'.��ɻ��t��F�kBQ+j�:����S�ܓf��672���:<s�a�w �M
w �v(J�F.f�՘W���u�b� ˃���X�Yw��@����s�^i0�s-w�zW�%n�ؼ�i�
n���xڱ�[�>f\HH�ɭ�l��ܾ�N����GAƺҊ������[�����N���U1�<��� �ú��ցEg)Cn�_z@�Y�*�t�(�1��k�Ŗj�,�iU�Ve5S*.A-�<Zr�K�g�����%�75P��,x8�UscŜs���!Y�.�t�>>h�������#��e�[5�B���n&�Af��v�����ם�k�J�,�QL�#������vo���a��2v���ٮ��U�dΎ�Y�������6��튄Ta-�i��qp1�B��Îٶ0��g�v��h|쁵��n3�g6�M�n��D��e.�M��R��W-X���9�bh�g��q��֤
^.��p�tZN���ѹ's`�8V�69�'i���lM|�O5 a��N�\zbY��J%�E����Ѓrt9u+���:�O&���Ս�^"�Q�kF-
�Ui�#̕��cGt�+\)B��=�l�����h���Uqf��pα1\ќ���:��Ҵb��w��v[w�x�q�u�/���@ �V� �Z�-T�ж���_���	��	�3�:�I�+<�
#J�.�.1����`冲��c
`��~�;��<��q�t��ށO:�Ba�Bz�yb�X��9��Y�8��zS%���S��A�ērtE��G��2� �ϙ��_�[�e=2�1� yj)}��(宾ڦ
G���)�De�*�@Y�2X�����MjZcJ2F�"��,��q8�ͫ3E�w�;�s�M�x�wS�R��MA��<���w?w�Ι/��YJ�SK�i	_	�1�)ی�Ywo_J\�i�k��4L� h@���A*OA�V4�ͺ�!��0_��`�p4��Mv)6���"[s����A�am���F��6$MJ��n!�%�Fzp�t|[�7&�a�_p>��ϭ�/ҾO����,���x-������8�lo6��i����ckň/��4�w�	`�S�>�U>���Q�ȣ�8!����&"�`bC��q�x��1�Z�J��Ĕ҆ LA�����H*�h"�(��"(���y/}u���1��_��r�����:}w��?��>ɝ��{���^�M���0w��������y�rN2 <RJ%B�	(
$W��!  �~C��<����������˙�w���C��=�]�o|�}��=׋�E�u��^$��e@@�s�	���O@W���	��~��N����	�O�mawS� ȵ,ɵ���e��[�a�� !����h?0e�2|�Va��o�학Gл�	p+�?�Vl�#�^?��j�rr)�9�0jӗ��(W�I���y��槚I�eש͏�
�l�<���w��<9�T�<�d����s�&�#O1��|��ܪg\�q��͉]�B֫�塊Erm%V��ͩ�h��\��/)�r>��,�h������zڔ/u����<�+&���C�Üv`���q��n#�\F䎣n^ۺno_k�����pdsy�߀�`E�6Z>��_�Y�\�tm��*��D��@m�Ԃ[߹d����,|5���'�'!���u��3���7<����f�]�6��<��L&�P��-�F�!��UcYs��VP-0`�Sp�p���6����j�F�-���R�~yɁx��'����YSg�vcA�j�s��N�4���\
���R���x��F�SQ\�;B�^���[6�<uВ�F��*����,�o�L��&��ܻ�A�/.��r�we�E�Ħn����̼�S��0"5�nG1�K6�`��{#�2�l�^:ۉ�7�6�*��)��.ҳOi(�>Ie�u/7_�Uq�\8�.珁q.~Ԯ�	,J)@�aQF=5��1G���:�Ϻ�Ĺ�ۋ&ӵ����]�0)�Z^m4�/Zv�,�3��ny^�fD�`J�J����Z�l�1
��J�oJ&��
w�{h(�����,Yܘ>vZ�쿆�0����k��T�lY�e��>k���X�_B������
S]8�F�f�flFr]���y�!��䪋�XScf-ys� 8  ��x�۬������<��q��.��8����h�2�������|Y�a������i�~ǖ��Y^��E����zcϥp`'<��BaE&�D��<�f4S�yt�j�� ��[894���Z�d�k���V�P�M��E!8(7����%���?[���������Z/4�P���h��J�&����kf1�I���,ᘕ�n��]�
�f�TՉ��)x��rf�E�d�ޜ��e9�}���Qf�5����Y�)�eƕYtn6}h���Q���ט|��»@2��ty�\U��i��릮ad�]v����B��ĝ��d�L����\H��L��$�dP��$˷�z�ZybD�E.�*3
6�M����8�3��8|���ը&�z�;B ��Vi������s�q�v�v��؇`Ur*&��&&h�)%�)J"�� ���4R1P�ZLMP�A�Rb(X��)�j�]�k���D~W���W����}���&w��>g�jo&� G�
\�DH� *��Y�}���P����O�d���.��������T��#b90�$�ʴQO�!�\-9�\�S#"�9ZEW���5�V���d�e9��Z��9;�B�nͨ<�[T�e\)Bd)�Y��R���J��@X�(BZ-�}q����f����ۭPtjGJ��;����Fb�6��D�39*�FTi��,�YZ�r_9�f=���y{��}k�Zc����d5YMB�.nU��L��bf�I.��I��" D�W��{n����s��yQ�|;���ݩ)y.�Kch��C�vUI�Ǿ�ރ�잂�ow��A�ڞ�Bq]��+��.��ߺ�]�$O���͕�ס%���j�4���f���[�NB��Oa �5\�al�73�{{�Q)޼�]�>��~���ʗ~�� �V��j�eWшW��`�.L�9��-6�����N��f�fa�{��pQ���Y~[��1��Ų�����UT3v����Բ��55�r�'�rO=�2s;��W�x�\;����;G�K�F%��)'3,]X���~^���^����q)�����'L������77�!�"���xm�0�'$Q�>dK�v�rp��Vn5���r���V]��h-9e���l7�cI�
��-���(4Kq!�?7a�V�I�J�9����Q���V���|בэzWڑ�bƖ�*|��9#J�7W�[��m[̞�2���R��Sv8x�4/����eQXV����j��Ī����5]��) T��IOň2w�փ(�_�T�8�����X��`I�v'}�Y�F�1:����y���ݱK�e�]�`7*a,{��U.Y?7I�]'���-Wڰ�iY�`�~|��Ǜr�U?+�hn�Xv���%h�m����۴YwF�L���`�0a٭����!�V>i����۵���ZO��iB��q�*��U*zsFUиT(n�]g�ӄD�4r��7[ov�6�v�����7�_�3K���NV�Sn����|����1��w&���w�Ѧmx���Z+2{ؓp�
�.Ui���,��P�.il��yn&�,�̄�yN$�#S%l��%��n��]B��C5��v��0�R���;u�_6�y�����i��y��]�q�v�wEw�}�x�~ӻ��pB$ci�$�O?�q��Q�z`3���ϗ�*�H��;�=e0;҉gƘRE(r�JyE����+/�'�i�gY���VlNP��ya9�<��*�}b���]ٰ�QT�d�,*	Fx��#QeLQrh�BVxq�-�=�������������t�ֽ��s�\{nW֓���<�:�%��j��L��<�;o���v�u~_�V���i��:y�&�,:�bF�[�h����v��b&D!�2Y�
�U�TiU)9!"1���e:�\�>�	Ib���Y�
=�
�9y�>I��>�z�߫�0��}1O�)���"�>1���B$~ǗL� �~����b��U��Bj�jD|����[jUsW5s�YV��.��-�/�ȡ)(
ibĦ!h�
\eH�+*���}۰�O�}�Z`"*�������?{��_�����7��?��#����>S����_�G��3 G��tx/��߫/��#��4�M$�%���ܢ�Y���\���W/f	&�^Y�!��F�VZ������%�>�Qj`R�S]����D�$p��f�mvh�B�`��Ξ��j��XyfKYX|5���xE��XvX"9����J%AJ�!U8{�c2F���Zq*�)�m)V�̢&jP��V���%U�T9��F98b���d��P�tD�u�RF�+
��VErpOu0D��`�(�T��pn�PHn��2�v�
.�*L�L-*Pb�w(��P�W,��ى���]��L�C���$һ�5P����`�*����]��`��jC%JE��j�C2rI%W!R����l��Ҋ.ZCKܜ0ay�w��%�L�!��L�C*\-�)1�{"���t�0D(�m�Z����Ay W�����K���;>����[���;���;˛�-����)��E�����q�駧a�Wf` ����`r�=�<�h�U�a&������ߞ��� ��(���+��s�����禧�y�_  <��e���v�%�5z��<�s)��Ŏɵ;���EAq�@�=���E���rpl-�!M��#�{�%;��7��pVrA���-����V��1��T�)u����x�l�m|����Ú���p̶GƁ�!P�y�{$��ıjsCI*�4Ӝ/��~��bڧ�e��+"�ԡ�b�{���j/���sSYB�:ԺJX�\�e`���C<��>=X5��ËGZ{٦�ha,"�fx���yb
����ӂòr�?=�٫�~��b=-��ŉ�x���ʋߒ5�|Ċ�{�q����f5Q�[�R�*��F����Y��R��&��ml;�s�����n)B����)�*s�E����KM����˞����ҧ\uup��s'�@�������ɮ杅��b��ݕA�庮d[����]|d��	t_��v����p� N��]g6;��m,�tOojS�˗�dt�&83��p,�o�N���$:wL��o}�&�4���8���R�Ʒ'e-�Z����ª����Y���Op�j۶�_Ƕ M�&<�\�Sw鴛��6<C��%�0]0D�7�/{)�p��	�6h�>��Y(�J_F����ы2;*K@��n�^�6�c�oY�sBZ���1�wQ̿#4؞=p�@��nyN��I,�i"r�r�8��O"�پ�X2��\w�fLSdy�s$�6��\X'׭�16'���8ϱ��)҈�^�7d��wD�pJ���lViJ��Xƙ����q�<�f$�ckv�C�+|
ѧ�O�e<����M����)���`���Ln�q�3gH�Ow������z�;�S׾�1���c7�؎�^�I�oLz�Z��!��OR����]~V�pS���;�^�S':���;O-K���+����/5�%����Ҡ��t�n��z�ߕt}�PCՋ�����F-�<h$�"J4�݊w�D�;+C,K�>�����owf8^��f>��'ǽ3��?m�����{��Nw�r���O<���)Q�n��:i؎��;5Ǹ���4���;��'��}�E�t}��ԛ�=�]8�n�X���=uO^���[��}}�Z�����>�q�̴�����'T��h���ȣ��t���� Jc���
&j)h
h"ij��eV�d�mF�jF��:Z�#M[m�S-�-R�غ�����)���}O�����߃������޶l���?#���O�OO��{�H#��@>%(|�N ӨO��9-ù8�L%D�1E4MLU5%$%TE4M13[�6�gJIh�ZS#"J?�����ɜ�������{���v|�w����F����v>p@k�yf;�	_�d 	@� R.�Y�繉��?m۞k��.�m3�]���b:z���EB�n��ܽ�'i�KmV�+FL*ƞ*	q���J�` � � �ғ�&&�X#)��8.���x�vE�Y�&��>��j��ё2��WQ3,*�ַ��^�r�i���ek�0VĨ�U�%��A���#��M�R��U�-��9'_��E��W�fk��2J]�������r��(��vF�Wn�v�ۊ�J�D+�L��wLމ�-|����(W|�i,l��P��Ȏ���N���+���ᣆ�~��ǤE�Sc�ro�ż���Y�ܧBr��d�f�oņ�YJfd��S�vG R�|�����<P���h���d@��nK�y�����x)kQl-.�Ǐk�I�T�v/��xF���
�W�mUPe,۾��w]�K�H�&�`1�f�OU�Q4���eGqk�2d�����A��I�ܔ5�75%�ce�sCn��ӽ����ǒ�r���
N�d+�i��`��[2�߻aJd]�ISy�N�i��)�l�~S�N�8���I�Yqlc��i�͞=�+&)��8��Ж��(��An���
�����0rQe2�7I�u���$�d��óN�۱P�"�Ħ|'�Mt�ƾW(h�w�N�q^��Vj�6]�=��yQ$4Q4�:�Q�t2�n�ҁfk��L�1�y&��;�����i朾�c�e�J�5��m�V�-�]ۍCF�?-��N�'gӵY�Ku������m�/�%�a�F�++���A�:Ƅ����٧
ķ��@܊��â�}������nP)�׀kF�&��I;,ɵ.�g=����j��vjR6cT�0ޙ���c#�u����K���o܏�;�C߼������O�ϧ��ƾ���������{A!�dJ��o��?'���]y���o�����˃/�_��٦�#����;�~�3�l���#�>:q����-��OE��ה:nދ˭��;zx���A��D�x3OH�ִ����y�ջ���N��A+�C"�ӿ���w41۾�~;�5m�f��oDQ�ܽ���,�Wh��ўsm��NcTOQ�����z�v��^y;���M�9�X��>����w����Ke�꧙t��Ƒ���=�~�t�G1/ ��)i���(Tw5!���Jb��~W��>@�����s�y/E��������?]�z����������;����w���  6�S!�C�R��4cy���b��CF&��0�SV�-SFM�c)��yč�y�y��y�=g
kt�
Ҳ�B��\�����A��B�Q����EGuQrfOlL����Z1�!���7�f3WvJ������4h����R�N	C$���G���cEQP�օO(d�fei&�O54ra.i��� �Y�;�B@U�����5���;ww{�k���Fyj�x;$h�D"ziVA7F�HU��V�n���4_���������鯚<����qV:7|����N��A�7ڷ�S
�FҐ�+�-*"�Nf	&�,J��{���aOP��/�S;���1@����y�Y��|:�����W��{�{���Ȅ~y�����u����s�s�9w_�����1"��&J��R�..	�jM��VL�`!��1�����1HKb-8(0L�|'�Qs���74�����x��|�HL!ER����ȧV�W��u��[��CD`P)^J��$Ý�-�]<�	uvt�:j:PO%n�(�����J
��U�%E*PY$��R�MWvn��aZ$�i���TQJ)��=<���9!K6�ht�9(rg/.�EG(��T�
��ҫ�WO�l���sx_wѧ�o�+:<�?�����n�7�&Jcs{5\�bY��uk����W*
�����ؐ��%�<PZ�$X1jj�F.�9{d�S6���)ffM�E�99J���Q32�Ph��L�7�/EP�D�t$��<)<1+ݥ��!����#�S���Y\h�;��o�_���U��pȖEWt�U�<$LT�ښ\غ)�[*;���R�Y{��X!L��.��L�!�]���"���PD˝P��)�AXq��7�M���B���X&F��@f&�
� ��maQ^P斱p�Ɛ��h�t��eV,U5�WF���N�b�+M�Q(���J)�*iA	�k�n�G��� �}1������G��wD`좨��$�"���)e�*giR�F�%��c|0���^�_���+�U�ȌvF�H�����o)RWl��Qd�"Q!�s T�AU��,'-m36$ҢmH#[�R�$@j�2&��P�E"����TU i�H�$4�C���#4��j��������W�6x���x�<E��{;�|{Y���D�9�D�5���y4�οRfkUW6Be|M���P���kvPH�bj���p��$z�w�C=Zt����ZRԸU�{w�alU����Y*�2���@W`���E���4͒�W �)Tf�B�Y=���v��oo������B[�����p)�J��KK2��!���y�y+T"a
g�����B�@\�D�w��3�T�Sd�&xG4{6l
&��
�=����$��B+d��z�#�f`�J�E�F�K
Q�Ƀ��&)���HieE���J��)J#*�:1!�ɰgCW{����g)eޅBDB�EJ��.)ʙ�j���p�*��Y�=��[[k~r���+{�^��w���|Ң(���C=Ĩ%����.Z
�Uց\"��^Y�g�w�^�����|���S(*R֡�
��[y5�K������;�U,��mpqn�S""�8t�7�&�S[VSF$��X���'�2�yc��x�sRt�p��)�xw{�^��C���Q�d�������
���/V𦢨�<A���,BE�C-�Q1al�Zܫ+B��Dڂ��W�Uh�w0�dGV�j����(���r,��Μ���.�Y-���%��,�Q���ĵwN��L�9�=��p��|��tH��O$���9w:�xG�����}��lhHIir��,-���̊D78z*dVEPKݮ=\�!��Ի!kW���bo��"��Sٯd�D|󇤃�]�o�uI��[[`�ު܅�Ò�ʵCє-�+U�5*�gT�uK$A��b"Ē�*[��Wi;S��,+�A3��5��{���i{5���8��R�gD�v�Q)hL"^�^-	��P��¤=�4�ַA��-�!Z�$x|�Ȥ�����<��F��^�����*dn�J���:E�[�#ȕx��++d�@hlFa�ꈬ@��Kr �d�ȁ	ZY�c�g��11Prp�)M�����r��eFUSr!��L���H�ga�����L1M S�&��M 0� �QK��J�����3UAU�8�IGU'��#Cedk�pw4�.�(ܖ�#�T�ܠ�L�f%2�jw��&��S�
�h���p�lL�V����MN]�d��)\>�|[���g��,�O;�o����S�.�lΟ<�\��w�MFT,���&�TȠj"-R"[م�ŝ��,Q���U��DK�-ZJ`�QB�U;FS�ɽ�C$:���Y����f!��.�XZi��u��Ҕdh����W7i'D%bZK	6��v�I�&a�"�n-�h�[D������v���B�z�Ɍ���Z�;�s`��ܖ���T���UL�r��ٻ�xOG'���`��)�t*�L�Y۱�-Z��y%6�4p��IXL�J�I�
�gr	%7p�u2�hl�kU5H1����w}-��j%��)��*�O:��A.l��	�.�,�َ&mĕ�%B�)��E�h�{Vܞ��珓Ф�y��]4����w�_���tM�ڋ������btJ���,��5ݩ3SU�[�g3EZ�WT�S%%T�f�O��$W
S&���"-MR%�ì�AS�i5uVy�JvR���)7h�n�2�md�;$!��%ZJ��,�L�Ԍ�-$UL�N�"Τ�!����
�唚%����+˳;@Y�$l��gSn`�Э)�L隅�9�)Z�jX�"�nF�KX�`��K�n��X����hO��m[�y琧�]wJ�Ζ{��\�(_&�;�w}�us�_��E��DUr�n`���z0Ln�w,��$��DS��Wzj�X{�T�"��d�v��*Z�Q���Yլ�"��kWF��u�z[��64bP�I�e"�fi��T����"���u&�JmiW �J�AQ1�TM�Ӥ<у%-GLj��a,�\�m�%���A��<�:��'�v]�׽�d����I�3���Q	�36(Sh�%��� R�D�!�*�Ѫ�Gf�$�al�H���y�eV�p���)�!��QB�2\̙��`鈮��쥮�<\P��hؤ2"����JAD�D��i��픨���3��J�7���_����	����"-�/����ݨ���^�bk�:w����[�Ѕb]ҽ�A5.e�D��j����wx�TEf�,����b�&NKD�m6��f�fܕ�մ����Q:�=C����e�R3%�C)g�v��hϕ�9�2R�y�/���Vb�6x�B�/�k��?|:[���g�+�t���V�39��KQ-t-�()+�FL��7�2ycT���0dZ0���L���ĚB�1[5M���i�!��P�!- �
Q�-��	D��r�qP�j%٦�M��JC�X����9�T/k���zBꦭ-�O^�Z�q��������`�y�����U�y��%-"8�j��%��Ζ���h�ou(��R��r��)���f)٢��Z��������|�.�{����z��`E�N�ea�!�<9A%H�%���U��glI͢�JU����h�6Xk��4/3�V!��BI�J4l2�+YS5�5��Zt���zrIT�������ܜ��ފJeh#	�t[@Tn����E	'A]e,�Z�%	��V�YTL�$Q�XgFeL��6b�yg�zup�
�I�����mV��.�2�i�`��,S�ɥ�v�l��Y�Z4t[�sfG$r䰪+�R�I[X��+CVI�'Y��0����f�d���`� �I��6IB�^]��)▍��6�l̾��w�'�׻�b����?����s��zKwfv{i�S4KʓYh��sKHg�GB��RGC��p��v�N�$�N�J;��[�S<Ӫ\S�2:��dUt��YY�Y�$�fJhkg�0��ؠ8�L�ɜU	&V��FBk�TxeV����Mt-iM�Q=��Z�Rce2x`���:C�3���W��������O<�W�{�.�U�}��e���嘗B���FJ|�3٩Zʽ"�5����(�fD���&5�Jý3Y<C-T�R�b�a�褎e�N����Z`�ڼ��^RV����|���!��5^&��Z(<�r���-�%V���$��=I�I��arqp�d
<�YA�`�e\��f��ѡ���\-v2��.�7�[�UGt�O2j�uN�4Tԫ9KFX���10D�0�Vt�4�U�m�gQ�wt�T%��	eRN�4nnU��@����<���=��U�x�&�4t��+6���ES`����tp��8G��뗐@��g��N�H��w'%-��-�ZRբ����ҝJ99��z3��qn�j�H$�U9�H7��6O"ޥ(�E�+� H$��N�̂�T��B�:*"�v"xP�k(F��5��v�+V��n�YcE|Y1ˠ��YѠ��S�\�D� ＞"R�=��z5f�{�=	"�"'���#�y�WB����䤦-�)������S+�e���-.�F.�%�c,p�kjP�-(CU�� �f�0ƕ6v얛����w�w�A����.=�h�3|�s؇�&�G�n�Y����\��7e`��RN��̔1��4���2QY������f�imW �����T�,"�R��P'���*�"N�'0�I����R�vf�΀��%ܖ������'pSJs��MU�W*��K��WVE6�f�.�.	�P�B]=�ZIM��Z����*U����R�c��ޜNZȘ���9`b$��J"A�Q����K�<�\�ܩ�LĲ�[�*ѓY�=3�2a&����h��х�ã͡�Y��=II�%"Κ�l��-J�ysC;�<����8�;�-~����7�&��eޑ�:6��O�s�HIx��><>�<W��'fw����>'�W������Uw�T�j��{ԳβE�K�#��w�\E#sWEA`�"�Y̩ю�����P���p�]>+�[�\�G���S>z̤��H�ҙ�B(���%J���j�m�W�nr����l����H������ Hl�	2�KKL�\lmYյ��m2�JčR�@#F%q+@��,�4S�1RS@R�Ҵ�HbV�1- @�"P�%%U��$�0�PX���ѵ`��$KJ�����`���mPbEP�5��-I[h�(V'�RV,@�J҅"��LBRP��\T�����mN`sQ��ٰ�X����������&H(,"����*d��LM�����ii�
v��6�hlM����iX���
��M��͛F���\�Ù
\E4�%	�q$GJ5\�̩l�����v+�M�+������zs���	ڷ�����~/��{_i��9��k���qv#k�x8�#��'��X�� W|p�~o�����sWxwo�\P�&��d�Q�%s���E�����_{���r�׊��l�n���8� @>��ŗ�z��g�f�f���~O��-H�я	�$�W��r"p�]g�֖�Â��J)�Bvruqʊ.\��d��[	��h��@��\cC��v3���AxA�s�>��1}1sƋ�e�-�n%�X%?Xס� 4��FY"�;��{/9��\�δ�(�{(�z����ƊÆX�=)�&]gS-�.+#|��¶��7�������������ẑWp=��^�~��Z9�>�㸳	`�K�ZF��_z�7&e�E|��K�i�E��\p�r�p���!gV�1(}����&���E�������YN�3L�a�1zba�a�mg�Xs�s��Y��WN��7F���ZJ�&���OJf�}�+O^ȝ$y�E{»~� �֋��؂�u �:�Ƀ>�M`�Q�F����!��\��π���.*n�Rl�	3�%O!���'Tǡ�n+��à��B�X��NTn&Έ��͠����2H�M���x��m9��|�ƍ�(�0g�6iT�[Uͺ⛏Q[��-�r�`t�绱Q(ѰPك���ڦ���\��=�Ƕ-����u���ٖS]�qJc77驇��q����K�8q�79���������}��uÓOq��<7�ze�+�Gu��ʛ&�8sCi/=�Wm���ŧ��\��*�*�����lzv�z�F��4I�r;���v�7�KJ4����3���rs���p�"E�Q���p��3X�H�Ӻ�(;�ndy� ��t���:T�'�Y^��&xg�y�5�Ӷ���k��Sc�9��<�뜉9��6��g��κ~��/�����,�Nھ�<�oxgmL���!���8�S'Q��uo.�G����w^VϪ��E��_����'��w��M���|T�:q��qƻΜ�M_>h�ʚ�7��cJ7����N}z�Θ#���U�2��l(n�eTPx6�u[N!'����������`)?����̪�S]C�E���­(R�	N$rj�(HĮo��o���}Wl�k�l��6�E����ٽό�;�7�+����� PS�̣��o1�?-�e�qv��>'���=4���Mb <��M�������>>?4Y^c�-Q�}���{.���Z�7��aD` �j<���2|<Ӊ	�9�K]�-���'>e�*_3�x��m��I��2�٘1�S���� W����JuCZ���!{&}c�wa2��3��gv���U��q-�3����������ݍi�Ot�w�wZ�՗B���sl��Tܯ��30ww0��Zu9����U@���G;uꅷ
��0��f�ߜ�͞�Kޛ)8�t\z�qgM�V�n�qן)Zv(-�"�U�#�堭�Μ9��������i�:S�l�#|ܢ@z�^�����&N����Z�0-x��Ox�%�rq�mK>ƊTQܷ���d���R����G�L��!]�˚�E�>~l�$�mM�'�{m���0{�sb^�hd��ş)�ȣ�,��'���y�7>|�(�K��J�LZӄ~���L���5�K�d�n�Tm[vj3�fK
�n����!��\�Ve���o��RN�:R�8�1i��\'ywu%s\ɟ��u,�"���H�?�-�y>WJz�:�{�9�<��iܜd�Mɞ�!li�V�r��vp��Y��Tc�Yz�?�8eY�hQ��S|\uNQ1(j�KWTf*냔�p\܌VD��Ǝ<�p�b��B�N���W����a��jϭ�n�b�MR6ϕ���c5�`e3��t��f��ʫT?[����h�5��F��l���8˒��nnd߄��¥���j��M�Vַ5��R؛k!D�Z09�R�OY%x�0%m%�ښ�.f�hՅ�Q޻��E?6�d	�9̺Oר�^Z�LřB�`�P�TW���0�Y�z��uT�|w���Z��G�@ �1���������(c)	g�p����L��U��'Ȫ�]�Y���H��ܿ&���2Z�.�ٹ�]b.��Z���@�N�dP�>��7G�.�Hi[@gC#O9>���B�>��2�|wL��9��szC�t﫻�~Zg$}���m��}O��E������V2K���p}pT3�YC�Ȧ4�6���Dra5LAP$L��l񅤨d&�h��|���'���o��������/������d�\?�|>��z����zX���}'es���;��  �$<ޑj��i�����|����ϖ|����1���=�����}������㼮�Ru�G�{C������&C"*�����,!�x9\�ׇ�=�A��4���KK?w���	O=>�:i�E�}�0)��<����F��щP�j��͸��u�k�Ʈ��W����؏���Ί�I;�sny���[O$2$�W^<���9 R�t�q���4G�ɯCd�|}�!���```��Z���澝�x�bЈ�����Q&E�YV����W����̶�G��_'���`������}���N����7ٽ���߇��@�&T8!�?�b������Oܹ��v�ei15Z�0��e 		���q��.[,�+�gόc��Ɩ�[J��쑗���+�h�a>Fp�mJzj��s1��}��MDp%�*�N��6�aW�8I�e(�"�*L MF���)��0��a� � ?`1�r`I�}���]QFtA�#�\T�`0�"�"Ck�����O���q���K�{�����_���~;�{��������j������C�v>��m轞" ��s�y �FA*�
9�
l��}��z=2��G��C�z���y�6��~|���p�׹v�
�1����s��{�~s�4��[�����{�ٞ��q3��Pǔ<��|�l�,a9��|����@�s>�3 � ,�c�N8�H�brT�C�LDP vi�BR$q���v��s;o��=��_�'7��o��w[��o��k�ޫĈ @��!ޅ�c>y0SW�>�`OQ��(�QKY$J�a�ɽ�w�@?�L��S�����yb/	��ьb0N3�'u��O��k�Ku��w��=CD$;��h�5���FJ
^y@� ��y���ahz�d��y��� �_^I'��ӽe
ߋ���أ╯�;��<_��{�I�?�=�:ӡb 0:M�A7.4@-握�Ֆ���{�*&�m�(bDQs�M$eh��WL80f	܋�Z��;��'��Vw��:	ώp9�</Ӟ��p�Jf�	�_+�<�x:|%f�X�6� �������_�ߑ��=��}v�C�	�K�����q70IV���}n�#þyÂRi�`�����@D�2��������� k���"|��˜�4��l8}}��C�F�łD��l�A�����p��ܟf|{��>�F��d����aCc�]��d�����y�s����
���T`
X�	��� p[E�wN�p��&"�@\�Q bc~���Y�V2,Q,S�1!��9��H�e�'.e}�w)� �F����̚������dO���zG�eg�����a�AA�{i�g �9��:��<�
���J�B�bC�I���Cl�� V0����.�H0&5!�	;(@/($�	U����blK�V�C��,�@��C�����}�}
N������C��J<�>|�!�����M�OS����x3�d N��a�%�蹘-a�P,Ũ� U��;��s݋a��i����gև�`w!��s�ސ� ��iId=��$�=�~c��Nz����_4��~>4r�Yl����|��lL�'6ot�Cl>>��w�>O���C�l�Yl���I��,�@P��ar!8�!��0��[��oS����-������*�O���;��[&U�Cs1��M���LɩF*�ܘ����f,�|����-�OF��{f�3L��C3�5Fm>��}Ҋ��S\.�'�wU�S#X���MF\�\UQykτ~���(ϫ1����Պ���Q?A�4{F�^��f�&��Q�n,yxbP�Rݛ�M�������UX̏����b+8Z�-�=cO�]7sEt��N��,Y�,��ĩ���U�p��L���kiOͽ�"<��L�������P���'ן+�}�\Ju)�-[K��=S���A9�̜N'-�'���3����+ǜ�ͫ���#�O)�Tu��dSt�iC}s�;ؖDꉦQ�Y��8)4�y{�TY¿g�>�}��cJ]���/��έ�ofCv��3tu��^pr<ґ��9m��o9�������������=����YN���ۛh��/X��VmvSA*���,fq��91m�K]��m�
���m�Zۉ��.Ӈ�ƿsM:^�{oM�M:n���Q�M�ɩJ.�sN/
#ӧN�q�- Oz�-i��zs�IH�۠�(�v�R
T���!
HH�Eeх�ʽ87�9ʈ���n��ܤ��F������VE���y����
��s��������~�>�����6��ۻ�5�2��"8�J��r���
fP�E+�i�K����4.V)�U��(�	k$�冄���\�th�;�{jx>O�y�""�E��XfRӦ	�@���(���(�w�JD�:f�I���;ߟ;��4��7n�����e85�V,Pà�)
��$�
h���D(x�xQA��9wsq��+6�w���ΕJ�w0����0�"�y� �z8�F:*:{y�q��Ny��Ӫ�T:^��(a�p=	`ѻ�\�w	E���<�r<Jwf`m�i�Eւ_~(�����p�Dj$�wgG7�C8�!� �\(8��B>�B�;W�Ü`�Wr`�<���(T���Χ�����N#�8|d٣���۳�J':a|9��3)Pm�����O^A�i�f�m���@z�8id��'�ħ ��m��W��P��0C�������<�5���-P�	��!�%8�hˌ_�y�o;@� ��Aws4]� 1�E�\��=w���"��M�?��O��{ϐ���s���h`@�Q�ѡ�p���}�yF���Z ���^:y���&	�	�i]��ŪLxm�SEo�4�#  ���p!�s�г�M�K@���`�	�&C� @�;WȀ3���V�)�{��;��a���p��8"��
Ä
�889��g	�z&	N y|=��#G�eA��٠��w�9�����0�9�Y��a�	�a��' ���g�V;F*�%B��m:F${c��2��4T- VM��]��sa���ɕ$����4;D��HLo0��̠�w����V��=�.$�-�`�
&`d@:���
Æ��e7$`h�)�i噑W� �hx��L"+wj��i�����9���:�Q]�r�5�L��� 7>X.��� $�E�p5�� �S˜�Q�� �L<�������7�9=�,���J$M��y��<c8(x��Y&"���9��Gvf0�I��{�����P�3���$Z7@��4ܹ^��p@#}�ә�� �h�g �lgK�������9��8?���9�N���t�s	fZ�3/{ѣ77	�!"<g�Šy��;s3�Y4ۙ� e����Ϟ����G�	���o�&C3��|�Cd32ME�Y16d����3'-�C�9&�����{��̰���&F��	��V͝aÜ�.��d:��O]4��<ݐȆ���}��'R�Y��������{s�h�ݚN��M2K�[4�Lw��7���ǜ����&�p0�L� e�z/2�P�=�I�,
<��9&P�p�D��qU���dѐ���
5����;M@8osY4��u��1
����s��Zؼ��b*!Ӕ2�d�A=��J��st�3M�Ӝ�1��gw5X�+�R+E濃�J)��J��s�TUM�NY�6��b��Z��k��_���8�����:�s(qH��������Ƙ#��q��M�.�u<��yE�4c�t�GGN��c�(�.�mMw5�h����P�ϸJ�ke���a��*�X��Uf
�o}rsx�&�ܕ�i�Fw�8qx����MU|�m3y���1U�ϧ3Ķ·.�.ٯ��U77U�<�Dݵ(e9�QTWoO\�m�p�C�8�+1*ee�s��崻����L�q�-]<��py8P����<���Q�4�M���t�����J4���n�t��I��g�Gsbw���ʧwv�'yN��0G&p�Ü*�i�0V.K��E�&��Wh�̜LU��ūJ�]2�C;��8w�����n�>w�خj�Fh�<�wV�0��h�8�D�pޜ/(����ʾ����*�\Q1���ߍ�g���M\��(�D�5pUp�
8w��m�6�����Si��53�<6Oc�."+�
_���i��ߺ��Q����<�ĵ���gV�ߎnQt
���$t�ގ�ސ�!Ojlpv�|��	�m���^g��|�k��f�<�ݔ�;_]�:�A���ӄ�uډ(�%b�M�M��5+�K����ޅR��}�fy�������͜��k�ᐯ>�qWQ���ާ����}~���ʾ�󽣠�w;恢��(�d0��� �$�ty�4Twh�����<G	Q��iMh[��o7W�����5��o%(����q���Uxi�wYj�^t�X���
M��4D�H_w� |�s��/���t��G��Wz{��!�sE�I<�d�.JE5Qtf���/�Nl�D�>o⏮�w����Η�׽Fҟ����þP�8�ǣw*�qA�	@��n*�F\�Ӂ�JF�=l�ְ��ü-��FR8q��ѹVbD��_�y�u���瞂�˔Q����pI�fm��~Ny�E	�xY�(~sN���O������]��5M�ӳ��Q���S��s9�]�ݻ�!Ϙ�0^+��Q�G|7xVf𛲑�\���4� �#{���t\�0� �&A�v�e����'(S����`I��H}�F!� Je�iRjFE�����I5(adVP�D��{.e�35�6���.��QJݑ'�}&�x�����<k�j؟����_������y�O��j}�*�12h�����#'pC�M%+IIHP5A��hC��'O��T�Jĥ!C� ����)@o��M�*l�$����0�Y��9�/��o��w/��ͩ�7�g�k�f�g�]���_;��^��e�u���k�mku�}���'��G��H���I�{��A���4��� ��;O��.Χ$*i��T�d������_k���7��?����H~�����P��ڸ�_��tսw���'z~7���?��>b�D����T{q��G�6̈w�k�.C�G�V�ҹ\��,	��{uj=x&��qj�1g�_5#:���F�\M����(���`�Sk3�#?\ɤ`��W��e�R��Ԩ�x�J9��/��sV��P�`M��)�]�>�|O�"I�_#�}���?�#���~��~���!��'��-����FHw�}&�+�w���*�� �0��͍��?Q�Eׇ��E?���:]S��@�bI��^���T�eJ)JA�$2�$Λ�|Ӊ�S�{�T�TCXe:���D�Z���0ĔR/��QI�ʇ�s0��%����,\�$�@�ۆҝ��6�����*�	�K��~pa�ȁq9*�)�&�|U���������^د��~�d�ei_�>��=�G�|a��;�I��Ԩbo����&d�s��('�?S���Mɾ*Z�9�[S/��?gWINO��i�5ĕ@OM�<Q��3����\�Q϶�*�j���&�VJ�������9���i����O޺=04`˒����ܧ�'�5 Σ�&���s?+���y�u6� �Ў��>ϸgN�.�1\�� BG�{O��n��5����L(� �F2�,	� P-2�fP��%b�E�lD�R�Xr��b�m��JZ-V"["Q�H����Ԙ>�Em=T���%�P���81P��	
`�|_��-�\/��]��y-�ޒdij������]h�O\�;ޏ�vf 餈DO�?��~��x���C�?e�y�b�P��+�8��+�t/�>I�ؐ�}�����=Q��/50��B�"�M{Oy�0����eSד��I1����_���J�+_��J�m�+�h9<�0=�&��֢����ί������o��sm�	z�yG�~4��-秞����+�q=ѧ�����e����B�-��:Y\K��t;H~s�����3#��t�xq��=��y����,���=���������� �b��s���9�ދ��k�����w�ს{ïw6�z'-v��!��w����)���:+����5ԝs��?(��y����M����+��7޲�F"�ym��ꗩ�>$>;��#��&���/�����}�:_���,�#�z���{[���E����e�����3V��p#��D���=}����C�����tA��z�	���!�:��Y�|&������B�N�0�C�����S�(�����A�v3,e�y~w�s�{}߷Ϫ��!!$" PGβ��'���O������c\O:��`v_�ۺ�G�9������8�6 %��s+�	4g�M����-��;(\�sWx�!�?Y?��w��d�����yT�/��w��q��&q8$P�H�Y��t��9���
x��u:;*���Y%/��)~������{r�����]���_Q�C�:�7��Y�#ف��w������L=�D������]�!M���_6�7?�����G��,'�ﾷ��=>��hD)[ÞS��P�!��M0S1��Ƞwo���x����O�=�޻y�H;���O�亟&g�{ѣ9�6A�F���6a8ޚ*�ۙ'�X}���a3<�v�yd��h�_��|Wm�4��B%Q�g�=���H� � �ݻL2N�7�l�U������+�~���k�q�i�P��.���]v��w����޷�������l����`���<�`6c)�e/�r�2u���*hk'�#���z�d�}��;�<���d��\��x-w!#�`dG���]�u�n��|V�d�3l!��O�#�,j7�Т����5��IBELU�AtB�s��X��y������<��д�# �$4PPT��SAE4-��)�����AB�,������*(�����EQ����֥�ib2�U�
�Q`��h+�QT���\DIKJ��#T�R�4�BД�AB
D$K"DT��Đ�o�y���f�fF��)�E�	U�eY�����10Q�2��Kn��L�&P��G[0�9�5ijqI��2юe0-��I BB��[^�3-��r��sȫľ9S����~Ӳ<G2�I�|��eX�R�A�*|��q�͔���[�����mZX��f�u̺��ˊ�Z8fZQ����wpt�s7(��'ȒH�:�#"0$�Oi�"CJ�eg�TTE����b�XV����-�%�cr�V��9�CLV���� �0�VҌE������Tic�EQ*-���*�"��J��EJ�1EDRUSU1�iBHD��Hxt���V�6ؕ* [U��X#"�elKh�*�DXT��b$Z�EZTYUVDX���UaF�b�Zb����5DT�h#QJ�*�Z$*)V�aY-��ʁ$��K+
�
�ԩb�[iQJ�cl��,-R���
�e�Z���[e����m�Vՠ�%[%��V-*[jU�`�Eie�Z�F��acJJ�&,X�1���!]�K�)�M��C׶@>���5�3��"�����a�^�N��)m\��XL�1��p�.8�4b�֭y��Vs��dr��/.�ǜ1����mWYQrS\U�F�����m��1UkTV�*��\V궴a����������1CSL� ��Qƫ\���d��6���ڮ4cicZ�fX�]h��(]�k�%(�r�yN!�h��XB@�$$o%ڪV-�J��؈��TDѨ�{��C��H{@B�E�b ��լR�Ư�e2q+C,�Tt�^��HB�q��Rҥ�_�$B@0��I	�d�g���ҙ�[mJ[TQ���e�T�Pe��*�1���>O�:2����s�^ݤis�k�qg=�y��>��<|G�f{lĨnY�ȥ���'�>�*�o������}�sn1q�OS���`���ؤ������S�Í��s�6�Z��q�
�,^+=��ߝ����>���j{��T�N���Q�9��|���5�Y�&JZ�(ʛ���3r�Lh_��~�nS�Dyv����7J��:�ӦN����ҳxTS3:yz�<i��g�ge��g�G�>ϭp��{E��.�080�v����:����
�{w�X{�z���K��T�ٝ3�t����'�=g������?/<=�� �>_.ALyC���ϕ���zHf���!�0�0�g�˓����|���h�����߰�Bl���E��{�а�g�^�un0�L���H����>���9o�G|���	O��w�<�>��{!>2L�d�����釟O;=����=S��)����Haa��l��M�Y'�!Ld,#>w�hwޝ������ιΧ�|6`�4��w8�ޔ�+��ɮA!�O������KE����p�0�N�ܡY�i�C4X>����r!�� �|4o���2�`�
1�`O(���m�l�@��B�m�ف�u&Fқg���Ͷ�O������=l��̀ʞ|餉9��DL�<0lm6�������O�3SJ�39�]���t��H�������}9��W��$)����Ps�mZ����)ѣ�Y}:]�\2�!���A9O��I�g�y���i�L�J�g�nl�����CD��h��gL��F�P_L,3&R�r<e��W��8��9�Z��]gt�����:��ަ{R�|�4�����N�OI,^��xd��D�bQaB+k�� $B`v��Mܝ����La�LI���ã �Q���a�301�ʇ��c�zH,�￶g�v�6��{��0�z�d�n����}������ף�:|��`||��1���������Kf��x��F(G�hi���O>��A��(�N�|�ִE+*V�k
��}�2��-�7-�iU]�b�Ķ�\©\�����%+U���@���������g�;1-3n��]�H���L���i�!��`����\ա�j΁zG°jBpL6���9a�]�S:����T���dɳ5���t%P�M4&,LDE�y�Ҝ�򪊂����t�8 x-Gbp�9�t{-��Ux_^Օ���'��!Oofբ���ҥ��U�U-�1iTcU��������3���4J�4)J4)JҔ&,I�Nc�[C�MSj}����뚩���fvy���$��3]����4Q0Q5SM5	ݡZ���;F0V!� ٱf���G�p�\�46�j��6h[�C򺇢�޴����ٰ�xه��Nv4��C�{��˷�lB��( �(i]��V�h�SaT�}[���A���6��	�?}rs*��&�.��\��9eMAEPLQ%5HST�	ABSPUDSHSQ��������i�.�_��u+y�GQ����>�H�K͗F<�y?A�Ѫ(�P��C��dS��7]��j.)�̕{?�:��'o�0~�S�s�U�O��1_��RI���=T�_�a3�o_����=@�ԃ7/����ߧC�-4���Lz�̈́�t�P�@�m���FJ}�����H���=��w�����z�	!�0^o��+�oi��J�����+)�.X���I�쿷Y����4�>�>��$��EH�����m��Z'�8�E�V}}�Z��8TD�sm.gS
n���7o�����D�f9T��l�[l	��s��ﶱ�e`�!YR}���W�ɋJڛ!D�@O=hϫ[�lS����x԰�5��1�c���� BI: �%�X[����G�O�������:�q:�8ʏ����=�=>���T~���'c�޴sxoz|�U�'�?�I����<��w��`Z]h�i����ʨ��2{_����v)Sȣ�����_O��u�4}u�\/q�9��)�M'�^l��x
��d'{�>��t�r�cK������3�G��WpI>W���C��$'�#�5� \�@L��I��lԀ�2$��q���o��n�u�-�_�_�q�9䚫%g�j}'}>�}S�~c;��#�;_��sR�����U�S8���$)��(Ly�&���S�3!	����9���yUY���O����L�i�qޓ,�<�(ʫ�8L������Uپ����~��/��)�]<� ¾��5����E��:<��N����&�{�Oq���3�3C�v�I��1 ��?�a���D_P	"GE+�����_?�:+���y���u� ;����<��uQ_���!����C�߬o���s�'�?��}?�~�|&>љ�r�nx��c��ۃ�[^�e��<��	����8�U�#���f���x����F���_���
�B>�;��k��]�^)\�%O��.�SO>~ջ�X}�C�|��TFR羶*�d�i^�|ℸU#��d�VC�w�z��~��l�O���?�?�?����W��{�|M���M]���_��*����������N����_��>�+���ƿ������(;�]�E_����a$=�CK&O��Ѽ���%X�2{/3q��/��Y�
Z��?�ؽa��Y���W�x�i>2zÓ{�b�D�umV�����c���������=`|�>�
2˩^�?��']�/��>��w��{�M�����&���-N�g�N[c�e��?���g�W�/��?�/8��DM/��?�,i��f��T���T��:�f���p�h=u v�dP��~��%ֱ�g!uT���R:��U�ƿ���Ԕ����ͱ$�d�)UtY.�ln�ɔcg*���݇B$h׏��J��%�m	$s�*ykNyX �R���܎i�(u���)PN�|K0��B�E"�B&hx�g�%�nǁ��`i��x0/Y.Z�P`q�}Sm�X ��A�@Af_*�)��Nr\�2����E� �"J\a����ݽ�C��9����Y�W0u�;o?��K�gS��"�0�J��Ĕ���o>u�;\�w�poi 4��v����8G4ߌ�b��[�CR��sSf��6L��4�HCQP��EQF�m�~K%Y�5J�ے{`H3��Բh��e�(���U-���/��wL�T�*�aEU��2�V�EX�[2�Eb�VcV&Ң�R���98@6d��e�*0����c,�(��Ι�ߤ�t��#�}�-S��:dNsM��[&�fٹ5YC��=%Z��>��y	�ԺJ�Y�;���;��PQTET��EUQMSL�QQAI*i��J�U5L��Jp;]�:�*�,��:2s+���)�65�������K�l���;�i)dT�,F��}�a�&�<�(�jX#1E��2�Y]�Gm��q�B�7�O�	�*v�h���Fh����Ù3�+2
�Q�?�̪+e!������w������|N��MH���O1��5���H���AjQ|>�F"~񰄄�%v��?����\�"��J_��=�*E�ｪ=��Ї�$��;����;�Y^��ϼ�8��UU־F�,����
w�W����և��1��
�w���-�����T��/0�=�Q\���t�4��E3�S�MDBP�����G����l*�r����z�X��z���U�<�USGU&"�a�����ÁV��EQTQQ���UPDQ-*�U(�*H����E 7䪍�px�̻q�c���S�郴PsqB�g-� m��dk�F6�ß��>9ƨk��z�G��ؤ�8��Qwt�K����"�������^��W�����2�*Z"�ގ�� K+*��c���uWx8�!���xP���]] 1����K|O�UT���<�4Y����(�d�z
��<��Wwu>dU�GR�T������^4�̥�3�1�G���dj���e&$�4l�.Pb\݌7:�&s� ��G������a���v�_s�y釧��K�*U��^���~p���z_��^W�w���{Jz�E����O7�w^�#�L�i^7��v�Kߠ1Ǻ{��]?է�v�~�>�K>	�C��V�����ո��{����N�ҧ���������
O��)_ x#�{=KΥR�D��|��\�eJ�O�e�Q�{�6~A�A���\0��q�H�;91)T%&"�T��`'�|��鮀m$��RDU)@�2��HO�l��T��E�
_soFa޷,q�cLGo�~.@�p��q)��:��T&�;�[���������=|��6���?	����0�G��kR�"T�kR��bV�CF#�T���
KF'�
"�
DE�!b��l��Q�Q� �F�Eb0[JV-��kR�� ��[T3!KLTL,P�,�,*"��ЕPVAQQADUSQ5C`���tt�<��Y���ڠH�5% 43Q@4,��R�RU<��0�g�=/O8�]���\�^
|���'�y��n���"ط����k�>bJ^¥YW<�@|��� :|A�IKмc��;ObR�)>���=#�o�^��W�y,|���*{0�^�z�K|@�k��>!�1��E��9 u�)��E�������'�e�OC^�:��Fʫ�����j.�T6R߅?M^ʎթ�?sk�]�=8a�W�iW�����]=����>ڧ��w�<�C���j���㦎��<ô��i����[������s���gT�>y��yW�����ӎ����I�O�@ �R2i������A��""��q�&%4�/�?Ys�F{C�v!���**"����B�$��ԕtd��#R��ltY;Ӳ�m-j$覮���_�ҥ�WW[�"�J����$��w��91n�r��t��F�V���`3C���9�!Gv,����W�|i�$eu�ڛT8��yl#����w^�Em�:�Oë֒���{��sT��0�T��+��~�=E_:J~L��_C8��󨽵L�«Wͣ��/2�q�@�!�j+��[#�g�TW���]��;7��~׿���#b�g0s��h�X\��m.r��ޯ�t�0�O���m���)i�%`)F��hl����uJ�[����py�wJ���Wv{?Q�U�?� f�YǬ������$2�Ji"����Q̦G�_�;*p�Q�F���X���گs����S��_ߏ2*�S����.�tNNʕxu=��T��e�0�.@�j�d�J0��h���<�G}�K���y=�Ǐ)�>�܏��a���B��@v���5=#�K�ЋJ5,
-U������B> jU��z���'Z%y�ƞ�����ƃ�a��閫�dI��A��X	d!���ٛ/��'Φ�(�O[P���M��`=�`�$$�� }R���r�7��l.H�  >�����Y����]у��D�����s�O�&X�"Ol���g�?4{�x�}?�[�b��C	�0�ߗ;Ŀ9JL��!W*  �0���)�����>�ᇁ�>���op9F6o(*(vu�fUά9^܍�I^�dyn�)v�+����9�.��W��QU�V�*��k ��4�$�~��A��_��ݙ��
n��Z<�?����Z�zBg�韛�������kǞ��K�mVȨ�*�t�6a�;��Cp���~�g��۽��)��U�Ǡz݀8�7:toiL��A5�8P����=���ߥ_%%,�.���<(�����󓷿�*�����Ei}W`O�2uTYS�h�Ӈ�����ED_�<���%.K�IH��{�BΪ�S糆���>;0�-�+���a�(��7�FB�!� d&�,~A1�w[��H- |ߗ���nypS�W��2>���gqǅ��ހ��N����:���f��ʻ��{�q?1�X�YqZX�x�e�>��1�K���f�GhȣA�y\��O�������c��,�K ��^̏��b6h�1�O͛�Z���h�2V�?X��R^�(��p1���l"d��{�)�C%?�&���O�{���:��&[k�!�ы���da}'-�J&���O�/>0��<�=C��c�|7feܐ���]`̝��qfhS�V�˿�+���?���硵�q���A-�a<PG�f1�co"��BP�E�B$>9򘂊�?
=� s��p>]UEa�&M���=���fM-"�������0g�ў�0=�%�%5�Ƒ��=#�r����u�:�L�� �Az���_�䁻%MG.��DU�s��k�T\��~��7�Ƿ�� h!� 0�����Ps=WL��t���m_�?�����fI��	�BZ70��B?�����9�C)'�_7�ٺ�Wi�Zԯk+��8?�e|����}���!�����Ic�@vyRA�'���#P�V�_p2���z8�N��lRyXN3,��Xs��ٲ�Y^S��qFP����C�y2�����ɉ �����,�!��a~Q!����, d�7�d�PO����LV\�6gJ�����U�x���`tȰ��d�"m_}4.Z��d�����N��#lGɔ=A�V��RhHQO��z��1#�~�0��������7�zv����U�f` Q�8�+�+�z3{K�����K�������������{�H �#�������z�BO�����@�}�����l}Oy�x~�2 O��Op���w��ߏ"d>���~B~���R �%1kuge��Vg�e��/� s��$�����N�I���3W%��hҌ�8��Jm%�?��sg�+�99����g��<U�3�*("��)�B��*����qۘ�� �4aX�F���x�
{@�����0(�o� Ն�m>{@>����}(���\��?ϼy�G�2�CMQ��c�C���f����F�A��=#�9C��s�}��2�=z\�r<�������#�xc�<x���v�m��������a��2�� �>2�A�Hy|f�D�t�����>GX�������;�>{?聆{��?�2��>Nr�W�?�o�o��{��<S�%��?	���`&e"���(��>�ͦ��㢺'�ju�4�]I�O�A4�*m�_��,	~��J��$Fo�|(@���sfў�8�S'��іC�%A1&]�01�ސh�O���rf4)I_VĘ� TX]3������c�st9����?,�~����sy�g�fD��ش���<��{jW�ť�k�4/����n?����s��ع\�R�ҡ�2~��������g:m'�|w�1"���΄!��q��9�_��?�4;�h9�
f�JVdT��0����۩��|\ � |i�wg�����`]��E����K{�t#�]~��~��Ow�����d�y��1Rv�}���z>�������U�<��ʊѠ��yrs� 3���5^L�!����_l�C�N�����.�wg1���`�ZGQ�'�j����A�s��\���$�'�0��8��IIB��JT�(0��u�0��oDK�:�=�4fN ���H�.���G�>I��4#&�V�%�����~��'�J�]�M/F��_�6g�$;c��h�-�������_��udij�jj4�d��f�����{�0 �� �����?���,��~�<'��O�����6����'����T��'�i�?�M�Y���ؚb��+u%�O�~8�T�ɶ'V3ؤ�����v7��IM`��z7n}��Pģȓ���1*�{�-QW���*�l_�^LL}�2��n6�EgX����� 2�Af @�¿��e���o�����x{�h��x�~�mMN�W(�;k�k��Q>����^���]�m�wh)��ׄI�כFKxז��¡$q�X6����x1��>+�� ���;1۷��)�0�ON���N�;�3F��Z�x���`���3�f+.H�L�V��gD��}'�}��~�왾_�_�}�⏛L�[��;o�C�8t�}����#�9�di�U�l�H����ш�>o��p��]7�?�������!�J����_�^y���x��O�.�ʢ��y��x���,�Ŏx�\덡ϣHZ����Q'm@����|с��     D {��OU�t}?��S��Lx��z��/�S�Qe�T�:�/֩�g^��Q��6�~Z��'��G�m�������'�e/�[n�9����yq�5�D��I�Ǧw1�[���L�S�2��q埁�Y�v�ae�Yv\ �(&��u a3��EI�|��w�G~�>g��O��������Qk��t�b?���t?.�G��j~:������!߮z/�nU\c�/c�϶�<s��v��|&���S��k�ϔ��|~��+��`��=�~���O�饦Hj��Bu���6��O�~P�Ώ�Ҕ�WZ��q͡��1k�mw�}'�|	=�X�2��X�2���i����W�W����)��{�{���4��/�i�k�F�������,X50̦�&��I�-��Y���Z�Y���Wm6�)�6lF5L��D�Җ��yQ�l���~���C�$�I'�w5s�W��FҜ�n�uγ1��ޝs����������� ��~nĒ�$� '����R��f]Y%Sr��0���[2)RYɆ*r�����!2�f��&T�v`�ջ�����=gg�����Q�BHn�V�VF�M,�M2��4����)���NS�|���PnF��j�?�UV�H�&�'�57VH�;j��X=��*�#2���o)�DS=�A�}AH��d3k�͉-/;#K�����Ò�ФU[eh�ϩ������i�����z�-�4�9) c ~`,:P㏰�b��7>D��Ɵl/X�gѵXеH�����;�l�?��G�>R��\�I払��9�.9F�ϐ�㉰z��o�h�s�V���Ȍ��Ά䚮t�,?U�%��ƺ�-I�=x��mo��tZN�G�rے� (�����0�
c}G5�.��p�f栻���������~7�"g�zg�x��8��˩Cu#�.���?a��[~�2hiջ�aO����>��\����}y�n��P�^V%�}+�t=;u݁K��
�k�Kݳ'�5�X׻�}���.u�PEŮ�/j㴧f~����+�N��u�L�w:?Y�˿�{����e�� ����~?3�?��Q*�:>�������m��~A��;�|Qyx�����篒|�W���w����B��Z�>=�tm4��j��N�Zuظ^�cr����{y^v:m�//���t���a��ݶr�g����s��co?�^��^\�ϗ]6�F[�����xm����a_}�<c���-����?;��|��_��z�ʔ��3FmL�Lp�=��[v�L�H�~c�D\
��	 eH_<�T���X�hj��*`�J*"���*����(��a)(*�����!��g Bʒ�1h��b�4j5~UʸA��*6j)�(�c1��::#r�x��2���$B�T�1�_�T�S8�\�0�$����}u:��
�֚h�80%UQIY262�a�-��H*���A$���rH�c|��d�����HHQQ螼H�ڤ����tG�m�s鰹/�\z�c������N݌Bp��:��l�)���Ck���L"�*I�(�҅'�q���.�l>)m�t�I,�4���2M�ON����n��c*h�8�Z��>�����n���$���h�Im�KDYF�.bQ��-u�`�p 5��g��b f$R�@�lo7�-�79p��j"^v-c�Y҆��� Y�LY��Q�lTT��6a.X�Jڔ��U*��jP��q!p�A:R�� �Q�K���*J��P�$k��D�&� ��:Vh&t���!6�	|T)�yiӌ��pT5(}ȅOJ��P]VY|-y#}��B7�Fx�)#I=�YeU�5��X�8e�QT(����`I5EYfY�zΔ�'���6x�m�х	ހep��=B��y����H�&��$ct!��ՙ��*,�kMB���)��	�COL�2qŬĬ�p�B�G�<��`T�q WʞE��P� �q�g��x�m�ͯ�����A=z\��QZ�EU������Ֆk��ɋ�� R?Iz��,�-���(���"P��~���й��I#Жq�R�L�a��M�]*�bi�Y5:�F�JF�D*UN���12J�����)R�2ɕ�+nG]l�Q*��&b�e�d���'4��*�36�bQG�1I�
4qp�Ze���9�K'�芭��U�g�WLJ�S�*�Ұ���pSE)�T����{�
+�#�Fj��l���}��u�9G��D�!#�7J��eW�a)`lJ�$rS[��b'O5a*���A:���ۼ�9����׉!����~'u����c�vt ��@ѥESԙƞ��~6�=�$��$���u�b�������tj�Ul�r��n9�2���� �	_�3�`��f���8�ʭbO�[�I��K"�4K���Z��>n�P�f*�]��i�Th��q��1"����K�#&�a�V�Ez�YK�!l�ZP��=�F�Mw�n��Ye����4���ȦeC�PVu�E
��\=\uQ���Gant(.��1��ZK�J�-��0�hՕ��igK��O��-KMD�m�eD+��2�Ͳu�Rē���%�fK���Sh�D���F"Sid!��V&����N�K:�\x ��ԐG+9i:�';q�Y��6Ed�nv�����5w��&��[`>�@x��;�P2��U���CSTɉ�������%IHQ����E�J#n��1q�o�����Ί�J�I�p�Y��ɑ�gyS�M�*gn��N6\����W
%���Z�N�Q�I� ��"��ĕ�ܒL�Y�k��c=|��I�<�.�Y��ؒ8(x�dW��l�,�9��%��k4O2s
�����~̵ZƖ��'��1EZL�`���U���p����S��2�6�a�,2�2�8l7�f�t4�(f-S��G���-\kP]�Wc&��8�n�ͯJU�z`��-�9o1e�M@Y7�Ǧ�Ǿ?*�mKf�ı8E����aW�>���nZ^�U�$���Fz��>C2w[�6�}y"�&�X-��	��lI2���"͆u�׎q�;�B�ĒXM>V��s_8�D7V}�`�0 �}����R5LY0̋���겓b`ƚm�RR&]��q	r�r��Ϯ��b�uJry�Y,�4�#����L�4��(Llw�����ɍl؍��|��]��5�Bv��z]M�^���o��d�Z��I)��-�#�,.>�E�42���n�؈��u:aY.�)�����ޖ���9NP�81�V'�W%�i�{����G��Ȑuьh�Q��Ҍ
��j�����Ũ`Z�.UU��X!<��幕���
�n,��
`W�'«��VW�� ��a��c
E��r��qy3>�F��A�Znl�!|�1މ���xṍ�������,e0^R�B�f�x�m���i�=3�%���Y�[UR����eO�SL��,��-L��j`�����-�E.��N^k�B��a606%�'�+ɤ@y� D}"����Ur����P �G}� �x=�4�6���"lw�a$}J�����B��hUL{2%�{"�"�0��٭�b1u.�T�l:�9�-����簱'�>���CtZ��Ⱙ�SM�:�;T����1X/ϲUHQ0ͬ�6g_��I�c2�E���������2�YY�7������ �@��%4	�7�^-J��#����3׵剺����EB(�ׯ)��'ΞՑ,m�XHX2:��q.��Ê��~�N��!��@z�bFY����l��iĭh��b��O�i�qG�i�&z[��ȤV�C�H�x�� .��{9�+~ʢȔƄq��Y�ʶ޽�-��	Dg�E����q4`��#���UR��BG��񙲥���<�������!�-2r���҉�g.C�����;5a�)�޳Ä
2�f��tY(��vQ��Y�v��q�x�SVŔ�ԷhǞˢ��&:��c��8�Ł��*l�+���q5Q��pA3Br	�(�D���6nC�X��\�"�ơkl�M����d[M�M[&�m 6F�V�I�E΍��:-�qЖ�jU�ZUB��SBSIM(P� D��&B��W)UͰ6�˚S���`�j�q"&��i�\JV��9��ŵG1sR���T��b�U��sS��4#��q�9��3[)�[Et�\�)�-�����)ѓhW2Q���U�T��9�sI[*檍��0W0F���@�5Кt��1Jl��4�l4Nb9�6 �Bڂ�JllI��ke["�Q�6�eF�lک��2��6�jNeljVԭ�[m!���U�[[�+jJ�fȭ�[�[blY���b���iP)Ti��16�����a��6��Bll[9� ؉sT-�T� �W2����s"lj*�ImUV�Sb��I�Q\Ҝ���e�a�ŴI���`��j�5Q�����kj���-��J�)[B6�s"�X������I�t�Fʖª�6M	m�sK�HsJ��[�\Ҷ���"s��8�ڍ�Q&D�)�
(@��C)LBД��� �T	J4���"�h���V
�UF����X���DP���*��
E"I1D�ҥ	ASTQBQT�
�ҌDHSH��5T�P�P�M)M P�R��HHR�II�DBPTMD����"�dUPQ@P�����JB��(�
iB�������)Z�
�"�Z

TX��"��m��
��IPQUEP�AU�UT�j�����"�H���������BSDH�QH�)AMAM4�!TP�*P�?{�}/�xo+Ｖ�o⾧�~����������������|�U���?��Y����cxz�!�GY���?��N󴺯�����������������'[���I�u�?��_�������v����W����;�>c�>o��t��U���`4
HʡB�ERT�C0T�T�KIUAQ@P�P$A��SET�EED��CAIJR+B� �J��f�F�6F��m@�J�JB�R�$�&��j�����[@h��hiR�hX��̍���m6ڛ(�(�h�hZ��P�*Db����iQ���)��)*��
�b*�J@�iP��hiR��")
h)V�$&�[2��l�6�el�ڛEl�إ�%�&�lCm�U�E�#e+jT-���ʖfiJ[6U6Ql��h�"m�6l��m
4�RT�SH�P��kjS`�6Dl��$�*&�-�[U*6�%��Ԩl�dTl��ڢl�(؄����&ŰHڪ[6T����d�6Bl��ȦȔڦғj��TڥE��h
F���i�
JD��
�!)�( �� )b ��$���(Fb��f����*��)����(��hd���i�&�i
bbf)"(��$�(ZlA����FЛ�b��6�m���a[
ڳl��6J�F�[B؛�-�[J��H6�I�#i[Y�Ki�6��e[!��E2�/����It�����!��G$�*�@��������c�3��;�a�=*��z.����~�}��=?����tI
�GɃ�{O����}�>{�>��]��������/O�;O��^����2ھ7�s������o����������}'x��}8l�>,���߻�a������a�_��a1}�����W���Wt����/����~�Q/�|���Y�����;��#?��{�}o����k�y�����s�?������>���ο��������?'ր @�,��S���_�ʮ�՚�fRP��A�2DQL�DT�DDD�QEADDARUUTPCLT�DQ�M1T�L�P��Q4DQQRS3PD�	L��EQEI$DEM%T�Q3SUDELT1UPT�T�ET�E1MD5D�TMLE4�TATD�L�3ATMLUA,E%AEMECD$�A1Q4QU5ED�ULATU4�QUUT��TSTSE4�Q1AJTUED�E4�EQMR�ETLIUTI4̑D�@L�PQ51QUT�4QSU0�Q%A����SUAUALQP�1UIPRALQLDSL�Q-QUQTA���PQI�IIE5TUQ$T�1L�UDU5$E4QTQLE-EUEUMS$S�BDQL3EAUPCTE5�QSM4KED�Q$RL�2ESUTAPETRUUD�TLEQASD��TPDQDT���I%CL5TQ-U11S�THIQEDET���EQE0L�RLATSDLE�SEUAEETS1QUELLUUP2QDEKDEM10U$�T��EDII$EPԐML�PD�LD�UST�MQ0STTPP�D�5I��DA4�MML5H�DQSAPD�UP0M!��� �徯��_w�-�������~o��_�o��j;����?�o���ߓ���o���s�g�}��}��xO��~׈�7�Y�{�Aّ���g0v?���<��f�>����k�����������}�K���������L[<�k�{�+���������L>��~���u_������{>���?�}[�����?��O��{�`� }�d���}���
��!���_D/Qؕ�����)��/�?�g�LG��2��+������>!�!�H����"0����yϒ���Y���ɞ�~�˲���Z��������O�*��Tn��l^��5�8��{�_���w�w�c����r�xGN��"�8�_|�-Z%�Ng��v69�O�!��qD�j,�gl ��$f�t�ꔑ6�����ElAkiŨ�S��I��4��w#��ΒG��$��|�鸞�]7f�ꅃ͔���N�����,@^��Eԡ5'U�5�'Z�+*D��ݻ6c�T��juĂ�����5�+~��c��RL�Oj9�e�\t��x4�")��z��5TR��WD{�k(ޭQf��)��9�,F`�6c&)`��Rڲ=rC���ػ�y��f��m[,5fj��יbG"�#C)'�MY�標���v3��� D������ܵ	4�Ǝ7%m��h�[�|F�h�==�k͞��%zk�b���A�7T�̅�H�Z��.
'��^��N�+^h��!�/�Dt�Gk "D |�{Z��vR:���r���_�ȟ�0�� ~Y
����T��s�:�_��VKa1�,�Ć�,$����+��B{! u��|���$:�S\�I8���,�� {���vHE$\}0�`H����H{��ē��a�'XO-��XC�Ԃ���fv�Yם0����R��������hɯLdP�`k$�r�c$���9��3jמ�Y&��q���:�r� OԄ��`������x�L8��OO�"����C��!Y"��%LBy�����T��(�Դ�VWR
])4�Ҕ1����}8�B��)�� zF23N�d=2zN�u= k��ΰZLJ�AH�R�����;��j6�i�T�)Q6J��=���+��+�S�BsQ�)u�S�:�U]2
:b�C��Ḙ���RsP�1�T�&����U<tx�;h���zH�ɐ>'YY8��5!�d���@�����&$��L���Md��'yIR,�E�$�!N���
J�V�8��B�x��D�l��1�$��q
�q@� HO8��P�LHb� B�PP%b�BIyI1������k$1�$%�B�=01��xg�;�����^9�lM�4�*
~3)Q��@j$����Q@Q@Ĥ����1AY&SY����*�������������������������������������ė^>�s�kK��±�\�� � � ����<����� >B$�(-<�m @ 4 h$� � P
 (=d ��    �   � 2� 5.mE( �}�[
x�H� EI SQ�����A�`f��  �q�@�@��F��ˀ    �����   1�,�  #X     �  4;�� 6  �=`  �7�  }        (  E  "�
   �%�mg� �np  �;Lm7�}nJ�C��mkB�AZ �b�
  �� ��^Q� �� �0���B� �!P�V�8Xh�D=ټ�Ĕ�y��^z�������vt"�X��ABR]�*������ D6��>ݼ�` �a�� @.�  �h�z @  f�����  De�    � q@XX͈�@       �i�c@4b00�!�&4�������OB`Si�l�'�iOS=SO&$ީ�)�'�O@
���?J{�G�	���"m5 �)�i�  �Pz� �4 ~��S@ d   @  ��h�i�D�iST���&�����4�� �4�hɂ�d�� ��aL LL`M= ai��ɀ �D���5(?T�Fʃ�6���ѣ�@  � �h�   M@�4F@� �@`@ѡ�� ��@�&��?I�2���)�Sb��4���l��='���O(���F�ā驴�d����F�P��6�OS@h����I�z��d��!R!� @ ��hi�ѩ�4h 4M�Jx��4$�dƓM`L�M�@4�4`�iS�ɦL#&L$@���t�	���J���R���Ǿ�B�1���HL�,|5i-�i���gŠ��^n�BŭdPr �a�"J�Ŵh���L��)p_iۮeMZ&���q���綽��V9巯���RY*xA6�l�B!�
H"��M#.���	h�E���5Ƙ[fGS�"3�u��<zI�o��������~Q �!O܆��~(�Nɢ���W��B|G��92M�}��~~��T_@�P����FF���ѫC!YM��kj��Pz���r�{U��S�/��&l��+ǖ?@ 1�a�Q׺��=WN��]������ט���F��u,�3 *�K��G�ѝ�����"�b �e��6��B��Y����;���ȩO}TW���M���0�_�?/������h	��i߷%�m >�(h�
ӊ�֩iS�|c����<@|�-Z�K>r��_+�3f�L4�۳��;�/8�#�!� x`(��uP���ڹ=�^��� ~
~[�������ǖcd�����>A�1w��+���0�v��J��x�z��y$��dVE�FDq�{�<
Z��O��i����P�J�0��Qr1'$)	�VnU��O$m��q�l��wj"��:�N��H���:��̡�_�)�穑V��,�3>F��0��q��*�D�u*��"uH��Sr ���N��-�u:�HD�-"�,�Vy�Z4g������DTv�E	PWvk������L�|D���y��(�x����2�K� >LE� m��)�Q�I��C�Eb���)�`<��aKm��a��KeF]SJ��\�6�ˬ���ʡv�wz���D�{�h1����ɯ��yx�\>�t�N�'-���o � P�����SJNxǨl7Tڷ`�r?m|�"������~�n��zO�N0o!��eOv�a4�S����&��!\�"$b	/�VL�z(}D�[9��=�%8�/���q���A��8 �p�m��1��^�=��ǫ���yP�`!���M0j�]V)E��w�9���� � a�<�������d�����<�=<�
9�_���7�I��9x�B>����H4��{~�zKȯ������h��'��fG�"���×��kAmUc'�iR*����w�����~�^vq8���UU1��o�6t�M\5$:���^��Uhc ���m���lN���u��vA��% I�`n�!3D�@~�"�F�2j����tά�?y�'�q|z�����vM��T����X�_�<���y�":+C�|�j|����o������%7]<O��9��c�Đ�B9,͑�#O�&��v��p��Q�vf4Z5�	V˳�o������5����O�ۄ��^�`��ʟ囻U��/V4+~�p�YA���M�x� ^Ϝ�;ۀ�\�Pt���ϐ��]�����ؔ��\�D���Cx���m���Mh����!]4�Q\*$��j�q A�C/h�	�h���]�j� Aּ7察S�Î����s�C�=y�Ru']��Hp&y�:s:�ր���[s�s< *��5ͨΎ�(��	c�:��ׯ/
�"M�|���}:��:.Ǳ�Ȯ����Vt3C�	�A�?B�˿l�o�c\뾙���� >��;�y���<����S��\���kg\8�׉>Ν�Vѹ�ϝ�2D�bs���o�������$�~C��u�a� �4��&� ,��@�>h Y�EE�&w��K��k�����@�����ؾ�k�J�sa�~~{��/�������/�c�ܑ�!��F����}�t�.��0�ɃA�)=n㿻�;�)[=���G!�\nK F���]!�ao2:��n�RT�&W���zN��7K2�����rdH�ӇjV�|���	M��o^��6)S�v��vv�]�A,�0���B�'e�F,e��3���9����8�������ʠ[x�u��y���[q�wv��2�s]����]�%��U�
!�\8JM;v�`�"uF�>=6�h�-^��& l�����
������2�h���ò"z����˝�0�@��h�:�N��锠���[�b��_V);Ч��N�c�8r�� ����	�9���?�InX�.�&�(͹o�9�B���!B��&/�$�dć�:���T� i	�؉X�o#��cUIn�9�˪���H,��_����gL�N"{���6�`5�2�Y�L/
�p���p��pր���op�M�R.���`�^,W>S�������8�/(ܜ��x�N9Ǯ9��c\s���p7n���RXn��LB��T+�E�)U�6�-���ׅ���fەU�\���,Խ-�[�+���x�6δz�=(�×c�#vN8���Hv}����9}ӊ���xQ[q�7{��k1P�m�1�gy\�EM���PXE
��ĳW|�G\��*6�C�N\����C�ܖ�F�g�*rp���Ȅ�U�%��K��������!����v�Ф�TFwu���FZ��ŤEW^h��U(2k�u|�kl:�]��Ց�s����CBxy/X��4��-'�"�GD�'9pTxX��q�k��$��s<�m�7�f��?[\��Td��w�3\�>]_^[��n}F)ni�'��53x>���ygOH��/��w;t[ب!���5p�+ϕӥ?N����7J�����o��#���[n���Ϗ/�G_>7Cl���ߟ���9m�M�О<��I�
zݺs���ٿ�r�����&k l��1��6�(�z��kN6�5&�%��f�����1��z��p4>o�^����9���F ]wM�/f/�Z�nCc��������8v�˱*-�wut=��p��Һ𯰩k�+��B3�_�� ]h��u���%:3]���(�,�9Li�.�PV7&����shE��-������92�����ǁ�� ƴ=�k�t6�q��P��bx߾�� 0DJM�8�VR���8:Asf�+�U��!��!H�zw�������o������?����}<5�AP4ZZ�}a� ރ�ƥx-���Ѧi;��O;�ɥ(Ծ°����[g�p}�����ÿOe>O���%��ȨG��ѻ��'���)�o�|G��z����GK�9:���薏
Ģ��&���z+u�Z����7�J�L_!;+x��ymߟ�塯��O~p�ǻ�3����Oe�_7�s�����n�E��������5^�����K)�{��f�eAD��` 5��$�44� 	���^8�p��H�Q�� �P�*n�۞/��pI(0)$�,5�­d�3c6���mm��#�yoN�kJ"C<�'+ J�	a40�����~g��5gW��@K���!�u�7Cց ��X`�ܗ�ucY��덍�����=?E��VӮ�E���H��'ax��*�S�y˄"o��o�?4�!��dq����@����y}�;���=?��|͐?��(�<�`ATǛ�K���~���Z�~���4��Es�0��Ƣl��ť0n�[��RJ�&!�`�N�R�L#Zx����-��<�8�:9�zJ�C#�V�)AC����i���~Z�N�e��TQ�w}u3���Y�;�:b������iJ�����������Y�q��"�z�4�%��@����cG�]��1&�o�.u'�i/���.1�ѫ.���go��׼��(+��������Zy'��}11~������|7�w��m���N2�<�I�>�S��sT�||:Չ�O�ȟ,'�Y�'=PHX�}�)�y�Z'p������p�s˄<ѝ�d @�3�XΚ�rg�o�<�O^>M�8�
myȴ&�P2�6�ʩ> �|/���Jg9���8C��[��2!2��hM�ꍞ	��Z�t�K.Xؑ��؂�f��"��)���P0}x� '�+��)<����L#��=��x��"#pz� �1��E"�'�Z7D�XAT�%�t�X�!j��Ó���;�#i��#�Z]�[Ej`kL�ud�"&�2� .4�5qp�vC=!�T��}U�	PN��H]���B�����u#\KRB9T�L��8��>X\�Š:����S��7���lL)�8x��T�(]���tFމ͜Bt.mrjp�����Q:���@����ެf}�D�P�I2�t�PU�$���x�Ν�v��؝������Qi͂��k�:(iݝ��<'Y�=N��-�N.r����;��O<�n��v�N���E�=�%��@ay
D-���i���ڂ� ҂WF�EٴN17��r�J��V����yz���tQeCk�ud��t�,���$(x�|�4��s����R�����˭4�Ze�ս��J�!c��tJ���.n��&�X�J��x�%Ts��Eoۡ
u�`�J"������1�ӫ=9kj���P�f���@�TĒRK
��L�O���*�3q)���cfdm��lض���)b�b%�I�i
�(fZ �B%�JBHba=Gp�PP^��ϒКbei�4c �&��e��<̬jR�U�8������Ds ��Q��7��z��xji���BYYebQ�J,��X����L��Ũ5Z(ju��8m�Y�q�:-lw�jh�@�iP���D���[�wƍoQ����i�F8��ˇ���t�n;��!EhB
�&�����a�r}q�����{��{A����A�O3(��7�����b�Ԩ.�4\�U��ŕ����ML�yp8Y�ק������>ޟ��~PW��UP����'��,o4
����p;}Zy=G��J�� fpx?w�p�4��8V�Gh�m) �  D@�Ӊ��zg���K����~/��>+���������?w���}��}�Y�~ �����s^��w��ߢ\��G��c�q�;��}��uYx���hf�|]Gv~_�����ޟeDS��5�}��'Y��yO5��yh��ټ��ϋ�5v+��W�D��O������ �i��
p򥥷V������\�0��q����P������W����{�?ϗ�7��7��5[�7�2O����J�+�����P$y��9����C� \���~^]���I�[��>^C�~���}W�	p=���n_��vؿ�d�u]v�E�z}/�����r|�������}_AL~����G���K麝�}_���0ί��o������G���z?G4�����3u~�w}����y�n����v~������zܿ����ߗ?�6Zb���__��������W����?�j:�.��zO!�>���O#��>g�ν�d��z�A��{��H9w8W��>�G�;;����3��yc�1c�p C���d"��߷ݯ��=s��u�vԌ��˹P�$
�(4�Ux�/�����}����L��.hUdx[n~��Τ���{�+��q:6x[��Gc��_���ű� l �\~�U���+��	�o�|�a����vd�#�y�v�}��R �]t�(�ӧ�z�gK�����hr�?���C���� �hh�:s߫6K 	 � �(w)�����0G*'�$�S��	\����St/j�ҽ`)�0Jb,��n0�D(HDȬ�ជk�{�X @�A A �y�A� ~��^=Y"��"�@k��=~�c䚴O���]z�'CC_T� D�=7���);#�z��׺�M�i'�3  p}KU0c�y2�BW+�=���A�$_��#����9�>g����MI��p�g�ժ���Նʖ�QMN� @+!�IO�N�HԠs�����J�Ỉ ij���4a�R�yI&n'� !� @ n8���Ez�S7����/M�"�:@ m�]k\��ߜL�D��-���q��i�`X��0!��I�	m@o<�R�}��騨ZA�e	ȔmC�b8��z�-�rt�"LH�O���L�ǆġ  �` @�:p�r�*�):���Z<���Q�u 7K ��<l��cO�}p'�4��Z���kZ����<ǃ̿#�w��}��|�a��l���OL�D o��N��9��c���	@�t�I�K	e	�Նp!�0A�9����Z �3�Mֺ� ��}��և�CZ֘� �|
,�%��53 �� 6��`��D�hE�/�
��b ݏ�,;�hD�O(�Ƞ ��ܐɤ��Ȼ��CPE�Ib�4X�R 	&M<��Ou�j !  @2j����Ld궓��#��и�~�#dr�ƑN�  !� *C_5J���`�f�Y�Ц<o�<�A>,��!X�8��9_wBe���$�Q� �  @�����<�ט���M6�u�J�WvtڶLR3*,���2G�� ��ԓ�Q���Ns(O�Y~���C%��J�Y�	("��6�$PV�la��!�$i)m  @
Qq���t�8B,�]Jg N	;�Փ2�Au���#�yt��q�N�A @&�΅�D`��8O�q���Q]?�Ն�EpҘ�+� #��� �d� ��+bB��	D���ډ&*A�  ��; �dNr�i��\��՝ꜷ�\��F�2�`�o�� A X���Vk��Pui(8޵#�Ӊ'Q�N�A @zɘ��xn�� GX@��U� �I���������<b�U[   �9P=UF�Œ��\���-�x��9���=>�����x0xv���CZ֐h��h�JP�`I,�64�Y�ByM$@ue�Wb�Q� �Cܖ��!�\^5
|�{h�̋c�pjc0�  ,�rp�-��g%
X��{�sD�����	�JP�Ҁ������`\���"�  @�K3%=gR5���Nʑ��ĥt/s ��{R!:� `N܉):���1�HwLA+�i'ag�Vl�6�.��ry)����XwQoF:���8z��l��� @�`d�n�
20 	)��.���Ȥ�����\�,����6M��Ҳ]n��3�E�9qӞ  �@@s  3�A��}B@t��l:I����h�7���`��kL2I?
@@ Ә5�P�:�SI;�t�0@� ���V[�'K8���(��Ȼ�����	;3�GXi��| � �y��.Q�Zȼi]y�D�6� �� @-^��A�l1���LX�`� �L��Z����I����#�pѮP1.�Tk�ܪ�y�i��  ���,��qH�"H�7���u��C@B�>*|����   A� #�y�����Gb�@�("$���`�m�aY$�+P�@h8���5������  �&������7f����b��n����ڣ� ��)��(� 8,$�\� p��i�i���ʞ�Aap�BX�H  ��F��� p�T�S?[�M��DD�"p,xF�P������p@��0j��  ���c���2���������h��E��S�����E`���GZ�zXZ�S��I @�� =)1�W�G
�NJ���B8��N�a$���!ï{K?{i����l�I��VH� � |В�J� ��]�AV�P1�8��� M��S�J3i��*�d�k'����t�	 @&�C9��d E�z�R�ַ�aP�h�ށ���!DF>~v�.F�e�  �6�%la��E.t��YN��p:�L�y��ӑ� �B  'B��O�`��C�Nqe�����IUL�KKI0�-m�\���Pz`| � �)�a<|1X2�8�}=�ޓi�?W�kC��>"����H=HD��v��.`x  �����xq�!���:\PA��n�$��I�4�dU&� � �=�t8�v�⫤{(i�c%��X@I�
.N�  � A 	�6.��{��H�o��&:5K<�Uѷ�&���� �i�h%I+rĖ�	f|�  �53����gW��5��&"πmC���A  @Ci���m�������~�w���+�6T��g��^CZր[��G묿G�R��15��=����ھG��ڜߡ� B�*�a�o�+�H�uW�Q�c�Z�-  @���s�a|��JԃvR�'����4��#�If��7�6Y#�z �b,��  �.-e�CIp�ai\1�N|�V��&�
��@��l΀m�B��|�  D�QV�0�D0�]R�#�g�YH�D��X�ǆ��(�5��߀�BA ���kV��.Q�`�7��#$C;����l� � ��Ci�2�j�E
�f�́Q��,� !� �<����D"  0��"TY�\���6%íH���r�D �  k@hq�<�
o��9��n)�{fףƜgDU>���W��BI� ��=	M~��3B��=Q�v㔣���a5��G֡�λW�;���Z��A-�:�Ơ�]��~>pg��j��mdu���{eD����np��;y�;�H@�ƭ���>M�S�^�ȶ^5<�/���8}O��x t����<D����n՝���˹�S�1]��[�{%�mm/ZeUo\%z�^�W	��6ݵw4\�V��E���$� �ҘD��KC��My[�J��B
D-A�(bm�����[��𠊒�V���K/�xsè��_>\ޥ���-�iZ��F
�]�Ա�[J�����
�٭o�q���B�ډ֝�c	��m���+^�媞���8Q���z�˭Fz�����b�mZ�Dϵ��>M�w4��K[+���%����W7�:�z�_l�=i�v���S	iO"e�+[7)��R	�0,��{����V��P�UG�wR�ͬm���^�^�ޭ�ڪ���Sަ�L�Y�y�{<k���k\5'5F=g�W�J�
Sk��w�+|�=��J�z;/{��3z�PR�^�����lr�*=L�;֧��X"(Ŏ�|�⭶�Un���߄�I����ƍ��V�^�,��KO�39�Lz��T=�T�
�]��2[W���d�Æ�k�q�m��~{w)�Ki�,�b^�MuwQJ���j�sϸ�k��֝�g]L9�YK[GݸxF��FZ�����z��|�[3�5/j=����Y�U�-U-o�s�̺��ݲs�T�YY�[��{Ty}��J��l���*��=NשX�گ_m���Ҧm�{`�3ڞ���U)2��4E�T�J%-j*0����ek�iuǭuYP�[�0�A:��R����ە*s�Qw�~;�|�{�U�� �SI ��T+x	��-ĀS
��k/HI /���˽	�|���+�����T#;=Z�kV1k/_j#�y�x���j��X������`�2@�`�F�Lu�!Dj���[	�YH�,A�K�>7u��5�-74�[9Z��n,������G"���6�b��>&7���cj9���v��벣V���4�ܨ�nM�ͨ�ko�|���e��d�UgX5h�M�Ͻ��{���jX�	�͂���f�.����m|�Ԭ�R�,���om��.��7Ko�ݹ:�N�LݖsF_�ƈ�*ũy6[K���j�3*]eG���ڧ7�\�qu�T\3������}��3|-t���������֦�[�K�븗�xE��M�kk�:ힴ_{��~{y%)~R�M��SF֕}5u��X���N��磞"��Ƿi�5)@�@b�e$�@�D����jUj�MKSSL�LI�Y&&��2B0$�y75l��ӯi�zsy��J��/yU����T��y+>Z&���A+��ɣNFB$���]��V��d�
㬗:���0�V��������\i��y��{�Z�C8<�)�-Y�93��}�R�L��n�و%n=�T)��i���!�9ϱL.�ޯ�;�����ZP�浮�4�m[��_{}��yo9�_&�ԣN�uV�7��a������E+����s�m]o��d�l����iz�%l�g=��Z�z�kKK��bv��x�^J0�����f��cf��dXa��U�Vڵ�6;S�:�௚�����罪��f6�ږ���q��ޣv���9��c��Ԭ��q��b���b�(�(d��P�=�f����M�Ui���͙*[_%��QQ޹���Υ�i�l_���E^Oj"(�֥fL��U~Y�|ަp�Zd�4뱪S�ʞsq���ŋ��40�T`�y6J�Pm,��J�[Y�M���w�7���M[wu�j��\(��n����|���u���"�>q�T�-Z�QEo�u��J��^��K�+�ۜ�m������&����J�����L�%J��=��2[J���T����۔�/�eUS5F=����Qh׵��v+m���3��l�V��i���Sk����h����*ߚ]j��Z�l#�R����Vz�9ō�+_5��g�z2m��2���AS*5k栊݅֏6xxc�k-|���i��*����B����V���+W4�Q��r���S�Gf���dɨ�
��l@�I��%��-V��rpV�>��dȸ�U�6���޽2���M=��a���TE֕o��F[Q���-_]֢�2���u,��Nx|כ�[��+a�69�ד5�J���ڬ���-��e��Up�J��׊�ҩ�{���Q�S̯�|��Z�x��}s��Z�l�JjvJ�N]DZ�R�_0��y_!밣[w�c���շ"��PEsR�,hYj�j �Z�x�ا��u5(suN��Yy��6ɪ�\e�����mE���kv�dr*U�q<��%����h��Z �a���wn��Yb�<�b�f�[Vx�\>���Tm�X=�^�ib��P��s<���v�l�:�'���qOR��-��"V�z�d�Q�ǵ�*QTe��Y�Ҿ��ܙ��U;�|�n��.����´lk+چ��ni��jU�UV�-��i�e�ڂŪ��+&�:���O>�)�Q��]�bԗ�.OS��7��b�G�nE}}��ϒ���]p��"�S�{7�k)�q��^�O\��ۃ��6�;k*��m[sq��<Z�]z�4n�׵�R�f3b����8�//�گ=�̻e�����/7�ɐ�j�wNB����ݭ�U'��|�By�*F��@N,�O����X���c@
�w�����2���W�eݵ�����;Y��;�|� o���z��������cc��'������\O��p6����V�o�����u������n?�!D%���w�#84Ɨ�n_1-*�j'a�&gl�CΏ�������hZZ�(
�h�f����&(j���I�)���!���~8�Y�_w��8����'Z��q;�w��<�jċ`�������+c#ɚ,Z� �x;�HK��@K�)*Q�ʵ��Z�g��/���:>�J����:�(J��\��%�_y�R.��G"�	k� ?��f�$G��{��.<��1�2��m]\r�Ӎ����Kඛ	Η��}��+mi�ypc)xׅ�r�)�>ڙN�wc� �v�mm��J�R�==蠲���5B��SN=[>��8�8R�-�g�-���Կ3�*����j�Љ��y1�8���d�l�n���[�Ln-����2�3薲uTI��SHv|�'A����z�GQ%��!����VK�i�ɛ6p12�eeJ���3>Uc�	l�ɚY(�Eh�A�����J�֐*��#r�����=\@�Cu��c�ԷQ3>��Bj���\��B��>�������jt��]���FՀƬPG�v�Y��:L��j��$���!�Y�6��qr��>L8�)�&q���n�1:��g��Y��mY��ݽ�k6�S'L�(�[j�^ipM�e�-IJYM۷���1�7ӄ�e�VzZc�Q��.�iXd�A ��~�9�!;*�f�B�*b��i
��bb��
�����Ji��f۟���5SQ���B8�[C��9ͨ?]�ގ��!�L�|� �_��������e}�Q��/9�~��η�7���*����=�PI8~�����U��?�T�>1�#��>g�~�(���e/���|�h����GO�Q��{jJ��V��4�)�gu���G��,�%*w��ؤ��6,C�!4{��{�<����eGd�p��eeȢ�7k���\�L�岯��tY�몼�NH+���r;�%a+K�6�Z6�v�e��L�y,Y1-p��e:�e�^Y������oQda�Le���b��Ǉ�k��9���5m˥�OF���Im�W����e��-u
֞��T�,�K,��/.������O;��?
���tH.5	�������62Wy�>r�*0TB-�倥�恦���+����$u��Ť�IEgN1R���Xϳ��,/)�v�a����|��U��j��:��9�.aJ+bsr���4�4&G�a��i8$ʈ���ʔf��b{��P�e�q�
�t���������r�ҽ�&��0�F���B�d5m;9e�J��&��;Cϝ��c��MO?[ Z:��j�ؘH��:���4!�\����h8����hDL�Z�߮��Q:6�.E<�)�J�B$H�I����|�9ϻ^�UQ�
'��#��$�w9#塢s�ڌJ,)a}�m��6���B�@7�-��4�ME�ޔ'f��`ۍ��{��saR-��:�V�����Zi���\r��jE6��>̘*D\��<�vn0��\|QV޾�l�{򮨜r�+Y�X�d=$����1dHM��vF�(
��u�V���z%�V��ެl`�9���q�6�'�؄I?K�W]��,7V8@=�� �$�kUT��R���g�Ϣ���%�j�l"lH����|�����m��8����/��P�� ���KGo�%�U��"��֤4
���HU+CL��!EJR"�P��)H͛!��ڦ��Q��u�I�?�ZZ�b���K��������*�-]���r��ͮ��keֶ3tB� �
����@ݯ��=���wN��'T�őL,��%��.��!�q��j�:Q��h����m(�~s����\���;t���i�kn����^��>w|:*����N�ɣN2TZ60F�����(a\d��[%��Vϓ{.$���{K}�U|�k�7��O���ix�L�'L�.�@(��Yp	�Q׳��\�Z���vЎ�@W�(���ݛ촅͵ ���sH]ڮm��������J��C�*�z�٬^Cٞ0��u�Q\ǣ^�#b��J�Z*ey^�ΰ�<mxb��'L�Y|�z�i�C���ߏ/<N��z��K��!����`����%^�R���S�I=5^�,{3�OM!|��R���<�RW���/o��5����w�O=� �����m+��P�G���|����ؖ�ԥ�6��j'v�dԋc�T����;hZ�S9�e�w9*[I��߀��B9�Ю�Lh�%4	FZp�P����#��
���T�p[G5*�2m]��H������q?d���Pt��>�~z�n`]s	a W(LC\����~���h����=_��?��u�I�M~��fS����������v�xo�������}�~����_'��zE�����Q�@�����t��%9Q�>�̔_E*�1/�L���G�� WMVL"�-�Y8� O��cS�0x%T)?O�^��K����O�����:�]�䆭=ß�U��^�p�qyq<f�3�ܙh�purѵ�'��p�&Q��[l6��{>�2.
��[�8��A�q�+ԋ܈�!��}.�/����\�/����h���I���ftH?�u�k�l߬�fO�}��:�M����;����U[���k}����8FC�3��@},�63 ϯg������]���[��e��o\|%����O/y�����Ng��-|���l�&�\#{����㺬��m�����ગ���J��U%&5:�U&����9�ʊ��jŲ���ĥm���Lś2ULPSEIT�Bm!�a'�-"�r���+���N?6��'[h_3��݀VyP���g�
��C�,$��� V��Sk�^���w��#�u�)�� a}��jڣd�QM�j�i�&�-�6	�+j��6A��u���ƦM�_�ӎ!*	^��{�y$�Hv�Sb��m[-�HvҥsR���m�� VNBI_!�$��� �a!$>0$����!̄3:���q�)�jM� ��Ĝ�7[�M��ؕNeJ��9����l�u���v�Z�u����ߐsR+b�HU��R�6�\h*l���2l�~��̒I�>w�3�"�U��0maZ�9�o2@���nDwx��'ΤMO:?/�l���"]F�^�wb���[x�׮>R�I�l�,I��"�!��"����i�i�2�"��Bk7��k��.L �[��t��q7ZH,��J��YkZ2q�j���z@M�^�B�cH�25����)�k+�;�d�q^ջ�iY[64����T���W��|�QU�
��ɓͲ�Z��ɓ�tI���)�n�۲��O�.��S�<R��m��|k�/4��F{�
���>����b����[m�ޢǛ>9�W���)L�eq֮�v>l�L�cPNq����[W+��;;���Q�Q�����ni�U,��)�g�u:NԢ�Jb��P�eOM��:�g�&��:�B� �cf��H��Ď�Dq�@�/�~3��U�D�)�I����)����s_;5)��־h�=�s�+������}�F6��׎ ���p��NЈ����u9O:ߝyw޸{���-zQO�����aϩ����kb�C��=�7�>[����f��ΐ5���A��BG�N�_��wg�kE��TM�c���Q�R�'���u�q��!��mܵ��ͳ���Q'v�3��u��,u�=���(s�M�l�*�	1�AƆ��Au�b�8��t�-�d��Z-aB�;+:���:���Ge����O���*�j�d�u�-n��i�����'>f<�9�Lʠ�׳E����;�;����k�b��ob�u۰�/ι(�Nu��m�<��x�ʶ�����*�v��o���
�jeK���2���j,m���2籓#�jW^ג����-��ڜ�|>�!sA�6�u��Aa�/��Z��P[E���Y�NK�L�,-�Q\v��_��ju�T��lT���wm���J����qj*:JL���ֵ*�{�ԑ�$ᖝ�9��mJ�mM(�Î9!���(�*�'7k�����R#�Kh�-�v�c�5;�@����Y+ fIIP� s$�e��Ӷ�9�8�l���\��!a�r���<��j�S�F��اYv�׎]�߅�GZ��'YM����j�6Kb��`�AƲ���������M�j��a��HwGyE4EV�2I���4�[lj���l6�dk5cM���)Z
�,�T@���:����,=����cͧu��2`G��0�>w�Y�f�2�<��4�W,��'2_�|����>�!�ty>-m�
u��������j�9���͞���0�$@�~���?�}�� �� ��?x����(�����W��R^�?��~|�G���G���g.��BK���܁�<L�D��t�hnG�: h�����������k�7�u���k�>�̓�)d� 뀿��fߤ���ɷ*��l��~���%I6��CR�:�I���W�S�2�vg�r�8805�(1AE&[|elv����=�ݕ:*.h�U�j���Rl6��بͩ�mm�a����M�V���2! ��6��i�lA�U[H�H�I�PsG5Nil���lxxfo�f*��J�#mP�Pg��s?E�|��Lab���Y�h�����sU�R3U�F�F3B�SZ]G.j�ԟkC��8E���)a�����y%"v�N�Ī��	�B�A�A��9T�y*`��RHB� $1m	�(ڋ�]d�dF,PQ�hr�)

�a�N*�q��ܨ�����~������W�8O��������߽ȣ/�)��|ߐ���}0�+�g/��c��9QME�
r�@L�
0�$?Z�S��TA}l���e,�E-* �
����UTUF��TY$�A�PɘQ���G%s3"!��
(�R栱AXf��0�=/4A�EES�$&I!� ���"�Rd�EG�F�TA�*(���[X�ET�PDc��z�����=�_�m�o�����s]��y�n��7��zm���v=�������|���O�p�`�����Q A�~�`��&Cl�QB��ւ�sPDYYD�  � dB,d�]|׋]_+�m��=?�
���;�C��lu�^�������/T��c����m#0���@@@�@^ p R$��	�U-������9*�h�k��5z�ڈrUA�P�r,9?d��X!<�;dY���"բ�1U�m�#"��,V2�*�%DQH1�9>_����h��8�[��ҩ��\��_E=RN8>в�q�Bm��XI��:��Vg���V��i�����I�r����GT����:�d��S	N��Dv�(=��}��Y�3c�U��M�T"�Ԗ����x�mY�ů^�Lj-�+�.5N�0����(�r�߁��)�q9��67�e���C/��\xU�`�u2�я&��T3�Y��V�\\�70d��H<{G>k�TW�J۲�}t5ӱ��`T�P)T`Ɗ_��k�rU��[���o8	�f�����.-Z�P]�oq{p�/	[
N�c �r5U����2�(�|В�u�̥Z�#�ٔ"�7�,�y�i�^��L%�U�RU�9�Z��D�k6�$��$[�[�i���r�!G%�D�^l�hTFR/�*k_����]�w�VBx�e2���C���%4��s&�ktb���6�X�אEmӧ��S&�P�?@dr���5�cH7��N)���Tǭ}�u8֜�O�	���^�4���wOA�a�

�_6}t����J6�^�HއE��r�:�ot�Ջ�P�K$aiW�y�oD���:;��b�:l��Z0Z�\
�OB�>�f���HX�2$��|�\VAgA�p:��;)k�LP����%�	�|2"�.&�d7�%Ε��T� �g��6u2�^S��FU�ל��n�&�2噸��M��&OU�߬  ��  �ѐX@�ђO�@:��Tu
�9ؔK"1!U[J���k2TX�(HH�(���9;R��g5�'2�Kh$9�ra�
J�P��wX,��L��������YF���Z�Ub#-�FՁTdP�ȕ ��D"�VC��I���Y �@��<�hT�L(�����
�s�Ub��_��`��C21����2T�������'�^0E�U(�c֨�eh)Z�̩�� ,��" �z��asFj��6����ְR���+�v>+��h��W�m�;?+��O�⸋_��~�m��Ll��]O����'�����O���K�,�^j�=��zHL1ו�SE/t�LB�~ɎG4E	n�"Q������AϮ��}O�D~�����s����=r,�х"�n�vAV��^�f��p
�'���m��鍍?�����|�ͦ{ \A��+`��m�l󚥴��wjko����P_���Ha��/6|t��|�e=䈺���Z�j�fJP2^�Q2i�=Q�[��mE�{ �U�J�1n$�{�^��lMs�H�M�ed�e���D�PřF�A
uƔ�ra�9]A8 �R�IW���k��+)�G<�fE�B�Z3&�nm����h�����2�G�a��ҚXt߃V�fiH�
���E�Wȶ�Z+%��Z��� �ې���4ԸMD�) *�w�Ѐ�T�)ﮟ	��u><Fp��&��9o�tD�4�Ƭ���$zCE� ���|n��lwXp �@Dz�Q�2��:�%(�t�ab���29�IYU�+!P���d�� p@��u���(
�Um�)E��r9I?C��{?;�yii������Ɓ,Ab�@P̄9 èX�ʕ*F�Eb����@�2s2E���O0ɑ���* 1%:$֌�(vi��"uUE��d�H�����*�l	�V-�X���� R��P���Z����IPY�*d!��~|��Ȱ����L�>08�1Y
ØX��Hd��U (��!0�U��*I��2EY�����|Ȥ���>pO�< �(Q	#h�UeO�`H.�RԿ�VXe@P����D�HI� 4�!)X�jز Q�"�6�*H+qB���*�ʤV�1)@`)%H%�a"$��[ X��%`��VB�(��ZYajQT%B�%�ZQjQ
��+V���h�J�J6�����%Z�Z��[Y[��dڭ�D��j�cRƥ��R��m�Tm
҅���9���U�	�9�AfT������
��C�P"�BrX�-�������EX,>��H|B
�R,d��	*U��"t؊iP3�4��)=�B��*ş�I�g� 2
�QX,��$̨� y�EdP��(,y����4V�L�@�aCH��(�Z��
�D(��C�ʦp9��c!�(J�	�J���d���}Ab�0��mb����	m��(}&@��n�H||���������>$�"�� ��RA`K ���(�8lX�S��2�� O psU`�R(��U��PP�> HYڑb�eD�����E �R��)� 6��޲��`�)-����L *��XʒTDtfYB�E4)U5H�4i�b�r�hP���fE�� ��e���#*�� �*I'$
�D��3Qn��
�s,��lPAm�v�ߡ�K`l4tfy'�Ty���۱j:��L��`��" T�y��f049&��T��Ŋ"ĕ���f��<�@{ǔg!Y*B�a֨��iV1�m��ה]jsb3]�
�<�#!�T��@̣}�v�PX�����$(�\�RKh�)2NI�J�ch�2(��
�EQ`���5ά��l�+	��a1
�z��-J�@���)eJ�sXD�D��졥W9B(I�u�^a3�U�bŁR�����5��j���r[���X���Eu�l�� �S����Qm9�Y�PX�����A#Q�"���a�̟ӽcz�Gh��mRԛO��0m��id�i��m�m�m���2i���@RRJ3T�P���R��Y
�hJ���wn�䝻����NC��������=�d�~S�����������G��w�
�� r�Jr�y�0ϭ�^Y����}�돴�xn�ʯ�|�Prj��5�1j4�G�Y�'u��/M鳼���gsgt�]���.��;_��n�b7˽����1�(���������W��?����'����{T=��x>��q�� & �=��gw�������|W5�ɑ��g���u&4=�~���߿�������|�zr���L�W�N4~�� ���3�=�|o�b�7����<�0n��ʁ�[��2�W�� �.#�y0���ԓO�U��ԏNa[��[vBm�([l� �}���(�'�2��y.fL>�3�J�Y�nz�gF�Q������P'z�?�vj�'�ʐ�ZǨ�X�v8�����}<:g�U�Np���V��b�:�;�-:�~��Ɖ�f�x]���&��#~|��d]	*}�����Z���(��}�5�X���Kgs=�sғCۅ��v�y6>%d�t�p��I�o2�tK�l�?���XSխ]HU�Z��,\N��M�t��$���ʙ|�_(�ۅ;Ȗ>L��o��s�-h�[�R��6W ��U�S�n��!s.��z,3Q�^|��K�iE����Z5R[]\�|lt6�p(LڧU�\>�����A\�_-	5;]��svkV鱆��G.��܁<�37>"�>�$���c֓�%o.�.��ƞ�j��Tn�ʯ9w�-�1�»��nY��q478�s7��|�ժ�0��م;.���Z�T0d�UG�{�|�5r�U|�5Q���i{G�V���f}�nd�j��DF�4Uo�V�=6ɿ��f�f��lGE�R��� �\�cq�q���Bk�~���<��8r)�qB�9B��i�3�W��m����ք䉂���dp��Y�}n%qΣ������k8�a^��6��ʶ�&�-��V�=弧XA�n�o�2� ��@?�$�=w�������0#��?� ��=�C�b�Q�?�3�!�4;O���'�I����>:~��Z,��`�"�7};�ҋ�	3NiUϺ�q���
�
�-3��9���L�_��I8�D�nZ�g��}Ͻ1�|�KFn��� j"_�BzB��(�I�cIU�����,�R`c+|?��H��Z���Fi��e��jʨ�E!�"�lF[ �\�N�s�Hh�N3�>$�5)ah�3##
��i�2��9�I�^��g�(��>LJ�J���������{V=��"���`���E��tB�oZ��d�Y��<���tS��!PlZ% dPi�S���xlm&�33�:z׃���%����M9��q!3�à���%�ɗV��Ys�`�c�C�m�,���Up����~�ɧS�@r�����K�O�iU��x��Vh�}�A��rj�4m)����I�Z`ɦҁ�?�iۿ&t𙨠�9{2�d���zG�?a�?��<���O�i�.U�Xэ�8�;=X�ͪꈪB�����*�
*��"�*�("�����j�����&����&��&��((���"���"������b"��*�(Ji�
iZ[�X ŉ��"�(
@�A�i��*�
"�h�F��1b)�R
DHVJ�PE������)�P�f�ԧ ���e������~��3�J����>���U8��^l������|_���}e�G"I�˗8�m�u������=�4 �_~u�W�UE)����DZr�h�j
���4����]WCq9N�ܤ�l�D�d�MFj6��Y�P��-KAH�5V���i�,����d6_Ng5*s.4[)��S��KAUR@� �����Z��G��O���3�Y������,����7��X���q����{��8�-�_���Sf��� �� �&`�U�"攫�T��l�ت���hT�sE��2n�CF�9�jјA콿�����������ⅿ̊���a�Y��/�� ���^�6�_��T?t����f���\T����P�O���X�����Ң���?�H �9�	��]��u<tj�R�kI`N�YD"CE��c0#��R�L��J"BJoЦ6Kԥ��r��Qa�X��)d�w�ZC �bIgz\~;�\�_w�U8w��>d����p�q}<>�:��[%=��C.{���D��M�_�]�����~9[�}����7��'&�)����f�x�v�ڔ��t��M��B�5r��*͜ߍI�oudiʕ�y�L�O<\_��R�ȳ���z���-��f��f��қ/G��!�5�.�U�?6p錺vN:߼sj��k�M�/M��Ւ|�ŰM�+J<��}�����1��(�S����hm�`�I�ݭ%V<��$��.���N]�5�at��vu�&j�U'��3��0�tҏ5��s�҂�K�c� ۱�ccsfl8b����&Ei�土���Qd��~4�&{pR��R)���GB���§����nb���y8��κ�̼'�����UP,�8�k
�F���.�V��H�J��RLPt���#v5xD�:��4z6n��x����o�:����1�VR�����.�R�n����2`�1#�;R�F%Kv��w�J"�u�Ӫ>��N���i.�!�&K�GF��Y���F��⺾I1S,ѫ� Ŷ����Vױ�x%�>��oсTn���M��ˀmcͭl�c9X�f���;	ϵ����r|1�UQ�W-պ��bM�2�\-Oh�Rf4�  :�  "@��{�,��E�1�����?&�z��}��|���{6��q=/��߼���ؽ�~Sݻ�������|��he�i_�mt#j�i�%�IO�ε��P���?߈�6��
����~L��+�z����	jZt���<r�&8C�<�a4�jA��l#���4�UY� §��$�fT���$�U�L��<Fc5��L�E�<ۗ�Q��?�I5Kd���Դgx��a�Hy%N���k�$��=T���+#�`&R�񟙶F��:VMTYU&r��]ћ�ˁ��~61�A�A�I���5�fe�b�	�B�ِ�Cu����g�����P�Z�On��jy-�{��r�J�OG-6;��)��l']T�cW���T���سG��	�ؑB�d%�W��XzTιm/!. 5Bm	����g~	�$䳔��"�9�#d�|l��{��o��~;�����|�xXp�Q�k~��WMv�|Z{�P�]��\�l�`l�F�f�j�j���Q�

B i�bb
��(J�C�����JZ�)F�� �ja"3UUC�����}G�����p:���:>S��	���꺍�M�=��~���O��>��\�޼�3����4h���'�e�V�����K��2�4��20�<���;�)��ok�^��O�t~#V�,x���>�sk%{�S�i�d���=�k������
�*  D,�����/{��?����s���9�u]�c�����]���dC�]��b·���ĉ�������UHedWu�m\��.3��|�����&������"fDN�f,�
�ǘ-�x&n>$��l�t1��j��kmN�s�����ᆭ�Z౼�ޠ���:��L��UYD-�?I̭���n����2TT�Z> ����Q�X��7��g9�i�Z�V�ɍ�vu1��Á�S�.S�*����+JNq��j}���2�|{��?D�Ů*ţUZI�*v���>ܠ�\��>�iN�p�-�i��\��9\7�=�O/�#�~��CY��O�'�i�Tm��.�eh���t=;�5+���ۅ�;�r\Gw4_�sX�p2�����H�Ɯ�F�G ���'��D���=2��0;�ay��~�W��[^����dӋ��rϣG����g�^�l��N����p�`�!���]agB����9�IL�B�b�&���+V�2�;�q��(ǋN���4p�I�Ǵ��H�����#?,�K[.܆�9��U�E6c.M'���}���kZ�l59sr�<u��g������;v�]��Z֩����<\�)F^Ç[';��w�ɋW�k5٢"��إ�5�o/�:��j�9�yT(Ѡĸ#�b��Q�:oO<Ѧk|�WKy.���["yz_�X�����+��˞�l��ۆZUW�/B�U�k%X�Am��oB�2��9W^�s�*�΀d<�Lu^rڙ1MAXOR���n}kl����G�^
���㎔��!���Y;Z�țȒ�7�k-:��� "  � ����$�� �^K����+��o}oy__�i\;�= 1 HaȮ�5ϼ}׆sj)�;�)���ez��4�&���x��*����f�ڠ���8Q|�I��%������3�J�O=�1/�\���`4(�xŋ�^~��gؓݠX���HX��ȧ:)Slr���֦�XT��R�����bQ ��W�.�&��2z��D��i���!��/x�J�A��UF#���I�sL)�qaT�#+�(GD�⊂j�/��Tf����Y�*|��H�AkU=7c� A�ܶ/Z�ٴ������<�G:�m�����$4E��z�X��X	�V]A�{�*4�Ġ��)�M��}[�au��:U�4-�L�����Y�\7�1����U���ĥ�L��tq"���� 	 @F'@� ��m��/rh��B��$bi(
���"
�)�����"��H&
��B��R�%�m�6��qQ41#�
���_$�~���7���X�^��x?��|��콧/���}?o����/�����Exc�� ?w���# ��h �8�=���]��=xwݗ��n��.`���?VwJ)Sx�a ��Q�}�y�����#�$�\y�Zw�[��Ŀ��Mo�w�?�}Kۉ�5�x8�ni$px��s��a�r�v" �c�5�[�:��М�/68�����b޸������
�	��������{#�>e�wņ,�d<��K�l')9���{.��r�ݓ��,j�E��;�mJ�r876[�.�t�9Zhɰ���B���/�%��Jq�0O�|P�J6>��,Z0�U�%���'��
�17��÷˗יz����V=~N� R\؞�+�c��R"�r�4��.8��}�am(eHsl�u���h����f�a}xs;�̇#��Zve�w�r�P۷V~L��\S1e�	Y�st�o�"��͢�r��A91������}��͜����^>��vN\�͓�Q6����;���	��U�O2�	*b��)�+�ӟc������^i[T�:Q���s^~;I�Ѷ��b@Ζi�Ŭ�t0]m���B��l�E������Gu��w�������#&���Y�/�dj�E�3݀��·��N>"��~���1����N'��q�h�`��lѣ);z�gW�љ�ō�y<��t])K��Ǔ>i�c~KS��7t�z�eI���G�V���Pp�k���#3�:O�$�5'O+)i�Yq}�m���N�C��}a
I*���yS�PȲɲ��xnu�ۯw�J���N:K�==ml(~�'I:�N<���:��[T�lw:�]ī�zZh�WY�hh��$���a�]�~Oo�w~!���6�	$VS�#����q��#�8�\��p�/�x�YO0Y&��'��'���_|A�Qo��O�����*ɭ�d���ᐽ�es �Rx>!��~�$f�ؔU��V��&�1�6\-��&�i7<W�>F��������ģD�s�(�@�ՉyRMn2d���R�RmQ��J��n��ôa,T8�(���f���� X�,	X,��' �S�D���m��,����iO"�n��}��]�5��V�m������V��Cq�L.�[*w��P\ ���]<ǘ$G�yL��% EN5t$h��@�R(�,�e���a�<w�r#W#��i8I�QP8I RFJP"bib�j���>�
� ;�����P�@�-QTSH�*BP�1%5�n�@�B�@�(��iJB���H�@�h�	$��	4�UQULJDs�_]��9�������=����S�\�����?���Y��Brq��I�b.��#�$�6������q��S.��P���M\	L������T|�* aW�m���LjJ�&�VlWQrR"[�`��)H�Tj�z�WK�+9�4f�>avVY��mQؐ�̭��A5��*��H|"c��I��H�Xdb�L�{���yK���KR��d��x�\*���r�i%�![.�
�XLyL�T�Ǐ��0��l�2�ٲ�B�SO��㌳��[;�kBi���Ͱ`�2;�g���WA�9�GI������˹q�l3�*�=We��=ߙ�xzf��}��E�	�z��$T�@y"�'�_�Ka��Wr���>߸l���4�
���#G��#�4	���#�=n�� 15ߕ��
��Ǣ�%�/}��;�{E��2v)��w��k��5�Y&ӵ�7p��V���d��E��҂� �*M��U���:�-��E��na�Y�ڞn�Dyl��$i�i�o�OB��˲>��,�r�kKr�/�$z7؍��WR�$�[���'l�q��I�V1��E6-Dۉs��=�M�qj��K��;J��9��g���1�*vN9L��&��v�|4sP�f�:V�͗7PR�N|XX�͙����V�aBwa��S7=��ej�Y�<�	5�mٝ����_�����֙J�%��ӞFc�j��X���2�N�h沓�6m�#�u�ޘ7��cC��F���"�q`���x�mV�v��s��饏�ک5�e���	/�N�;�>�d�$!�,}�Q]���ǝ%d��Z[9���sm�9l�a��P� �'��)��]'F��O�ܲ'QcF��3-Яw���msG��;k�7E
K)�!��ٞ.R3�u˪�tp9�ũʜ�eU�]ٟGL�`���h,�8��]i���M�H~^�iͱ�e�F�7"�rs)�+�UoG-���?�C�h��W~L8n�>���ޜi�M�׃�&�cCM��J��6b�ҁ�5j܆���*���O��O3�{iIp~�*�Jb8�C28b���-�@ ��Ȕ!wU�߽����s�w�Ϧ�%�~w�$�T�(]2L)�D�2�#,��U3���A�y�`��v�0��(=��m�J����9� �"��J���^�+�)CD�L�~7������Ƿ��~�
����7�η�W�솯'�*�Ad�$c�"�dN,۬��	��EM�63P~��Z$�Պ�#�,Jō$�+V����$�Q8{��i)��8�<��8��%!�tr,���d��%�(��	�!�����8�+d��]G��m �e6���{��!I���LR"���	1W�<k�\q��w(]2{��M�	EE!K,�q��(�!@��Z�'6���Ű�3�cb)R�DHE����{��������k��:�_�k��N�M���׹a����������?%�<�@ c�!a��c��>�H��~�P�38�M�ka��idG�T\�Ʋ�4*`�ܚFtZ,��ŝRY�AYaR�-l=�RYV*īT�L����_�YҜ�j�F����̒�d�j���e%�6V	.�	�l�G���1R��E"4�](������L�s�g2���៥�6�y��V�(��Wi�E^M�h\LV�ukk�W�S�L��.fU�c	�*j��D�̒ӄ��4����ؒU���9��%���	�Oyo9L���[�hc�7O�#(b�ZX@�96a��Цz��wdG�4�]���Qo�J(E-*ty�"d��Yk�EƑ,�(�����o�M!�o:��م��܎�|�x�t��o�wo��{�>����T�]XP9?������5����A}���m��5�w���F�s���n�:��j�SϽ�=���`��*�v�}*H �RM
������H{�mc=~^�]����S������I�'��2�O�������T�I��C8��3?�5�	���<���[8-g0�X�A*̺40�A}_.*e�Zs^�B#]������2�2L�)9"$s�����h��e�������5rǕ�O��v��q�îJ��@���a��E�*�c9崭�X5{fP�ej��W�:�޾E?L�v�/��[��i�G�>��6*to�*l�����s�o�zڎwOݜ�I��p�\w���<�V��7/ʇ���̦�T�IţD��%U��`��:p�ѢdI�g=��aD���N��ę��.�T����a�\sms��QHk%�D�O���F�Y�X��i���\IUrHڰ:���uR�Hm����xtV\X\�}Nq������,z�=:b�nY��-X���qϗ{���tin��1O��k���M��C�y/K\�;�nݳ�f̫���S���]�)�Nm�ߥ��$㢀�Ҋ�@�8w�
X��N�6sB���}�U��
*N\������K���υK-x�룆Oq)���#lo5;w��L�a1+a�V-��^\���Be��(q�DS�|��[�OK��#�M�p�y�bW{��M�'�,��s)՚8
��7ޭy4��"tb��T����׏kK�'��X�h�{���l�vDĆ�S�/�����@5�J�[�*�_K&-��,�q\Yth��  �#�z�^��p�}���`OnJ]ʂ�;p%�C'�u�z���H �)�Q'�-/8���I�,�ey��p�a۪���͒ �'�h��f�|EO3`�d��h�r�\�La�)2p$3ID��3*pJA/!C�0�+F6�E%,@i�iRʲg@������{��)5��ey΁h�P~�N��ҩ�������;.�)y���=���'$��3	@��@��)�y㕹�9��p��PJu(n
����/?UV��߆�L:7n.��dw��;��sǏ������N�=���瀆�£��yf$$�>��xJ���()�bT b"%E�R-+�(bJ
�� "/�c�g�|ߏ�yA��������[���燫��+�4?��{��ٿ/������y`��0%�E&#��}��y�e!�9QL��LRD�MIT�EP�4TETEUUW& �	I@���A�|�ۻ�#�;���t��q޼'����&��{���H����g�-0� ����i��ٌ�\܅�]r*�gî>�?ȡ���_b�"�[]�QԴ��~3����Z�* @ ����oZ-g��v��G\�w�)i� <��}�x��,��N���7Lk3�u��3�kXB{aנ��M �^y$�t��ap���Ћ#t�$;�ٿ��y�c�ǩ|�ɤ�3�Xˬ{3H��&�z	Ť퐽����5�$4�Ji�Q���<��k���"J�:Mcq&�Y+i��m�����ۡ�l�_Sl�e����;Z��4���m8�L$�Sd��&����	��v�7�H�gV���Y��@���lz��aF��Ƕ1���#}�#^KP�B��kꔻ�.�ԏrL��WLG�\5����6���j-E��/n�Zµ4�ѷJ1��O9q!sx��e�(�u)+�v9�N�̦m�)Xg�[�G�3�e�8d8�\2��R�^mOk����3���Qzp4��{v�M��{+�������8�&^�g�8���h���Z(����vX�^��[���Ž�#����J��c�͂�w��,{1��(�w��˺��S�I[S�4^�[�0�b&s9�hv��_ns�nW,}��=��]��YZ�:W���3n��1g�YIa׼�Ӷ�SŶ�9�l�:�mྫྷ�Ssq&�KL����f��٣U���$v���X�a�x�{=s_���H�$��\M���j�ڱ�ạ�^�VmvA�,x�V\��b��fs��1R��������D8@�@ � � ��%��o%��_Z_k�ܞGd�Mc'�;�1��=�[פW����= u���}�s���$�=�_w�y�gS�S�3���{8����V(CUh����z*<Tj,#��]t�-�^)��]����$Z'��K�Y�$!3"��.C�Gp��V%x
MVݴ{��}����z���v'��M�n�ӿ�����|P�؞�W�����Z=���ov2��J#��+������o~���G��m���Zs�n5�<ΰ��?�,�� į�OQգJkl͙��I�3Z5�V����LD*'}�W�<���_+���͎�����E�<������q�C��o_��^���8�45�~?��S����'���o�Ki��/��
�&f5�f��4����������I
ރ���{S��8���.�mm7n�yCoJ`��UH�^��b>�@��*�dKRHY���V�(�f���A�l�+
���	5R�X�BZqpĦX����5�UI��/Qu8���E�'ym,^!��L��y\*e�$d�;*\����
��6��
Z��f�}�.b�T\0�sB���ԭ8c,�v��*���j1E��ʙB��мcV2�mR�u����:*��l�Rf�CED�ѡ)J�M.W�2��@��"��8�u����½��0�N;�d�J�0�{$��%�8ځJ��a�`mZ�R���KZ�:^@�$D�D�Càe�	E.�U!P%+[���Nl2��i̊9�^�!/
CS�.X��8�*DC1�,���3�p�,�"�)JIx�-q��B��)/j+����4_�9�OH]�צ�;6K���+"uE��9oAi�!�efEil��9�j�[�����b�26(+b\ܵ��͜�`�y�+�6K��dZ��m�'Jئ+.��5+R���.PȁeHYx�le!b��e�&�%�"b�"ܝd�99��dU�\Q��KGE|B�+:�M6af���,C�QR..	f��*,[�٢沖�#d��j6M�":	���K�[4�H�i����Q��ىE4�ɨL�!M�W��{k�J��w��K�62r�$(��X@�)�D�SNɡyO�^�K�Il���j�v."(|z���
��8�4�u8f�N�E�H/R�jVIӵC��&o)L=��|�|�hJ�f���b"o1)�Z��z�t�iO���Cd�ý�bba��EyK��Jd�7/V�rY"mR��Rr�
3�f�#��e�-�IB�א��L�,-d���`�)��c�C�<��Lɦ[&2�[U�ܛ��(�	Hj\�}"EQB΁KL�����2E��S����D8�CE�d����s
��)�H�8DMl����=4mR���8�S�Cӭ̈́i���dT�I�6mQ��{D1U���S!�V�-��t�onEc.���˗�P���ej����R��ѪDwi��M+90��iRE%�NCLZЩ�|an�p!���k���Y��VZ�\C"���Y\�zJ�A�-e�1Xڴ��ɼ�KdW�8q;�2"�,�([33.�b�x���Iw�Ɠ�pN�e*�ق��Dh��6�N���*Vg!�L㢖P�B�b���-"1����f�	h��rڵѠ�d8L|j���D䵵�%��(�t��0$Q����ޮ���*'!�wuh�(��0C0��Z2�s4�.,:�J{(��X�f�\XK.���^���&h-��\=�]܄�y��B�*���b�H��6�p�XU��
�+q,	�Ƅ���0>L+�B���S=�Z��AJ3-m�\���b�d�@i��I��*Rm�K3�P����1��e\�|b�!�-	D��70�sS�p��-V8�.rCL��Sv�mj��k Z�K�;��V4���(�S+��M�ic�L�%���Y^�3-��+VU[c�J$��+(���yypnr�<kTԯ
�Ua��1���*�[��B%�TK���!�^K��<%4�Ų�*1�Ed��Vd��6��U�UJƒ�*�Cd����(�-���M�Qsl�&�"�+<7���*�!�E�@�n����n���Ыt�r����<��E�pQU5U�����5�+�6��on���͌�Y�W&���0�>	�{X�m/WQw�����C"��P)���,U:�[$�[EH�G8Uj"p�%������2�.����]���Q�fU�]���"QB.SP�g4�Kh��=Eԉ{����P4���ˎ�f̘G�Q�fP�E$5�A��h�]�@���Q�0�D�v�"�#H�*�4FT�%"��ՙ��������)U7/�v����dFQ-yj*��!Z�֞��|1�&jQ�Z`�LS���e�5+��\YԹwt�M1�m*Au��S�j2��p逰4�Kbbʇ�	�$ίj�8��)����a2����g$]��%�TN��!,��x4ʘ����.Ե5�3c^��#^R��O�x(�+�>�[JEC�,�J�Đ�l���a����F^QU�1{4w����f2)�;�����
;=Z�U̼=�+X�0��UUL�a���]T��e�g���\IaT�Sr�Mq+\�"J��i�u�i[�rld��9�-�&��%,B��!�V3�!���JI���rRZ�S��ҷn.��.Z枔W	"�0��E2�N[����T�Ff(�MK�Z�H��^�1@���j����b��%%�V0�b�ȸ�r@6V)��F>1�+0���D�j�2f�P�\3��ˈT��8�"=b�>"0y�M0 ��qW+*���"���-$=�J��"!%NR��,���Z�(ܜ�����z�C��9E�ȵ3�%��J���WIk8�b�R�4���U�Ӗ.�ON�ĔB�3*ʻ7,n�@�-X�F=�ie&qI�\0��ܗ�U��v��#*�d�$�PMe��;D�18Ҩ��0����NA����-"�^"ë�{t�SE��<�aYj��w�h(�mfY��,+��A�ƼUe��)��� �:�ų.�^�س�����7�����{K�Y��&��)����3��%\^ib^Ҵ��¬���.�{$%	I�ꪭ[U3T]���v�BB�E!�S4$���v��`ȏ���5R1�M��F��^.7[��З��龱9H������£��^����e�����0�(�%�.��ik��j�%�"#]�[e�j�2��E%�`���^�'z������Y9�;=V'<ڎŴY8M3��2(qf���SX����wʖY-�IOh�KX�h�ejļ�X59H���k�x����;d��gc"��I�i4X�̑X�%ݓ%�`K�3��,2.���Z���YrJk�Fh��dK"�X�2�\LI���ђ���&�	�heA��s��3�>;�S�Y�rb�fx�GyR�+Y`*V-PE���KF�ґ8��&��ԣ��6��������g�;I�X��t,�^=�F�b���2в���T����B֟2b����#�}=C�a+i-�3�,�3�xZ����%-�q�!�*��Q����UE�Xb�%.R@��%-���:J9V�o-�d�t���K��nƁWJ�!�_)�d��KF��U�|���E��Z�.�X^u��F��)U9sI�C���CB�]�����ǆ|XrR�*�iRb��-P!T�K2Hl%֦-��c�6"+0���-�ЙU���w�wv!&P�f�z��T���i�Z�̜�ÐBM%˙\�J��8��!�%�-�v�W��l�0%�lv��VJ*@e������%TK�#E%���Uf6���&���L��'9+��)C=Fw}��0=�=�z�>��O��E�Q�twzò{Ja;�����*iS�b��8q�䙧..��E)�f�P��a��#�2Ж��{&�b.X4���2<�84�w�l����\q����¼Nf�)=�g|�����)��E{��-��׍�b�.+c*Z�v奥�X"�-ZPy�P��2^U�eM�ʊ�rL%TJ���i��\���Q.*�4���xɩ�&��d�-=+3E��T���jm�3bQI�W���ʩ�1���
*@qEi�f��A��!����d3	
2l�I�X��v�iv5wZ�_idF��I[S쁖�:�2��Q����/yR8��Zu�c���U�E��F��� ��YCq"eo(�BB[LȖ{E����XCeͥD��|�I���X��&N/��f�q��||�N�Auy���j�3�W$1�]�;���4(#A��*�0=�ٴJ�	Er)��"aB[�@�Y�#gxuɺ�����{M�R�A2�s��)�PXHQ���gb�"/�)���4©�[���*���%\����)H�v��-�1-�T:d.��Xě���1��.Ѫ*2re.Yҩ� v�*���$b�&:BڹyH��-v���ZE���LX0-NJe��FD�^-�[�,4�JLI�ũr�X�T�HvVHR��(��ɶ��S�V,�@dej%�)���n]�(m(�8%T�J�g�bC�V�-7��K��Xȥ�($�4-țVL��h�Y^�(E�2��d
�5%��0�ȷyr�+0�=Z=d��L�2ҶeXAhK�k�R��c�6ƈ�.���N*f2�V�ma�!
-
T+oN���pmZV��º��;�TYdTj�|�AO��gD�P��z���J��K˜[u�jQ$T<����A���U���%��9��wx������|t4��*��N�-K��d��e�d���-Z�(�� ������\4���$�L������Qc-̻�(��j��e<��M�d����rR��,�9V�g+C�C�L�b���&A˔V�z���!T�y�!�%���*Y$��E��UI�L���4����S*#�^bU��]Ȃ���&%�C]M�(�FeZ�.)j
Z�e�gRI��y��Q7d(�[W��k�i5&�SD�1�&!�F�%�V�5���ا3j�4sF�j�9�s��T ��
+J��,HT�P����B�
V�lml[�jmff�ڣ���l6������H��P�T�ńD�0�""q�MT�4�b�����$J�E!@��-KHQ��%HVE�aUc[��46����s6'0bZR 1�\U������T�eAJ�HV#+�)J�(ċH�E��s6�-��ch65W2q�sI����[�� $  �Y�;��=#���/�0fy�p�?(��C��<�#�o��=&��U�� C���Q=7����%+vv�B[�OYpgn�mڡ�����l�r"q�����,��t��zB"����LF��`@xT���7���'D@+P��{�cFL+F]�7nɛ��Ik�1��U�+s��}�y�Q��J�,L��ܥ���"�͈շ�9p�[;����9,�w$��c��|�� �;?N��=��F��|���SV�ئ��v9�Y�Pd��5�����T4V�#q�=D�%,n��7�!��{-�k�k�l�k�Q�s�:m�,g�/!����GmnW�7RQbh�\9(��J�N��`я��[zm]�Np���D�n�����_Z��(iy�,早�M���CY8�QZ�w%Ƚ�-_S�Jݏ凊F�dI]8�Q�6l�����ɋ����βTp�k�c�݉����׷'*��kɃ�7��J���o�£x�M
.��p��w�A}V���9��].��Vk~�1����.g�����[})�c|UG|Nٻ�'��V��_0�6kIS1Jo2hAZŋ��I�Y�p��s�Xm�N�QW�������PVYJ�AE�VZ������̔M��y��Kk��2g���r��L��ޓ ��,��ˁ	�/R��cM�%�c�e���.$��� l�I�D�u�6ů:���s;+Q
�b΄v��3rss	�6a�=<����I:�v=�g�.�?�=p�5�r��O���g~�u'U �,h"���@u��`_\����6n�������K9�D{��bK8��1%��~d����̵�����c�yGXᓿӯ�������� �@��8D��
�'ǿ*�N�fU��ÒO���3���)��W_�Yq�s��}g�P�p�A��%"�A�)ec
4n���qߥ����%B'~����FdJp�����wU�yrq�����잆e���= ?��GC�kZ�}���F��eW6�B��H��
eE~'s�w���o��;�~��|�x��o��7�� � ��`D��d
~����&��%�ty0hzh����/0V/1�����aT|��������F3(y�o��i�>�K��E-k��5k��:Y�ߚ&xF/A�~<JA s��i�?+)t��
+�q��Փ�~�2�Rj��{�I%��v:�"ya��g���Ӿ���+'s�z62����=��Q؝���݇��ӗ�3�Ӣ�sno:Y�3f�e�K�e'\lO閍XsQ�Kc���:UɃ�vSf�ǈħ�#�6���wd��H`���"��}�\�����бLm^n�J\ou7ޱam�Ptgr���{>e%��.vܖm��L'v�e����튊�����ph��@Ms�H�j���mo;�鉛�A*�x�EjPݼ�S"���Y���{j����OC�f�7��\�e�BK�*3gӐ�GZ��Y��g�/��˞6ƂZ��a$m��y�ݰ"�����p��v�*�8kϧj·l&�L�6B���3n�����Ne\��Y����m&R0h������_�c#�_:V-3J�a�jک'|�_�p�m�[���47fY0�#�W'���].��3׿D�&<����R�6ay�Zv#��J�URM��,�+H�ؖIN��-En��P��.�r���ǫ���2p㖷+�F�KͯH%�
6e1�yj���.�x�4�z��(Z���{;q��f���陦�Y��]��J��\>���e���qjR�����8�g��� o,��S%�?���������8
T�ޏlS���>�S���<�䒰���z�����qlv�ǚL��W����/4:����D�4�DdV����좒e>������[�>����|l?=�??�矠�\q�ǆ����9yR�凶Z���_.��p�<�g�ϕ�b�$�|[�%�+Q'�LL;Cyy��/q��˝%R�I�r�5��R�l��ߟ}���S-�n^]��Ƭ�գV��ck,��0wAF0{r}�(� 9��+����	QR��w�x�����������5�~��s_�����<�������~��v|���',���KJ)2LDTLIMh"}����~���gc�>��NR��ak�1S�4v��c���~�}������5�u���f����]1;�Z�X;�>}s]��/k�>����o2����b��f3�6�'�׷Y��S|X����ֵ��O�5Q�&�����j����1��GU��~�zO��:?�����}���~s������ؼ���|wn�8�����ԥ�_��١ڬX0�a������jZ �@�k�������C7�_C�-(E���T�� I�!h8? ���N���`|�����(0�C�ؗH��	O`�ۉ�8	s��ei��ӳ������v�����&&��Wl���/Fq���)�t���
�������Y��~����W깮/���~_�������b��*�� ���� ��&@?#����ܹa��~|�a� >w��~�����0>ITQ���ș��	/��	��S#z���h�4����BHGfx����ՠ~���2��L &I��m�{�#�~��q������_?��>��w�{O%��7O�>O��>'K�������'�}7A�#�Z��Q���r'��:-\>��<7�ce�vn�v\6�c=:2���*���M~O�~%
����I$7����ҿ������d�A�^��OH�/HgY��g�th]�#�]�c�� ְ��ܹ3.G7�C��?��܉�jJ�(�q�j�D�@���ѝ	q%�J�.�8A���(L������
 >�N$�A~��@����]@g�h�-��#���(	�G��a��APB��r����Y�|�6����Q�/@��l$(|
���-���\	.3�	m����Dk{Q��ᤝh� �BP<��l�|C�? �p�7/Н6�h���@V��������
����<$c "��i�̑"h@RWX�C�I��H4J5LR�1&h�@롮��F�X`�v%�ј��A;�lP��Kg#HѸ<�ͨi��X�ε����-��Ѡ�4m8���$=���@N� ���;�@6�06�>H���_ ���� ��P� ��YH�!�;�9��i�*'��<��ɿ>
ì�C��@�`-�Q&B�Q$����]>g4,�����(� ���{�Ǔc�=I��֔��E 93�\P���=s�q1#��~/�hH" �؇�v��+���:�	�ݵ8h
�F���ˍ{?=G1��x$��*�ﾳ� �h�g���3�q� s��s�tpx� ��}�G곙>�}�|NO�/�S�D��-��j e�jƃ�d�"W �����{�`0YHYO�'�}��Xá�<���#��|:�g��37� ���~���D�O���~�	Y8��`~���6�0�����x�ۨ�(���V��k��bx�=���	�BQ
��*��%T�넇?��{�	�Z�2�g�)�+�=�SQg��#*Y�c�7��Î3"!�$��(8%�)$ +����c$�?����������O_�9x�x�υg��ޡ�wP��!��~��; �_n��lQ��w}OX�6s�Z@�(	 ��pM��A�{ǽ�Od��CM�y�<�h����p�%b ���G!������ra$E����!��y�n }u�J"��&b���J�D$��	O0K<�����B$�ōa�x��$��8��0�D�;��H5������a_(�"#)�F"{[�˽��w����|���d�9�SΞ۞�r^v��Pߴ6��>XH���	%�L�]&P�Iq�Z�[�y���H� 0I_����@w���H��:p&ILY��͵�`��DW<#֞>�n���^�
�}���sR	I	�`&�V�졈؂�p�!��,T�	��6�D�<�3WO�y�A�<H�p� �	%��E�wyP��Cۡ�E0D0�d�4�^�N�̑���-�(����D% �e���H%�y�2�;�� ��O$' ($rm�8G4p��#�2c���!ՅR�ރ4�������L�.	{�8H�O;G7�
[brL��A����Q��]AVz���L�E"s�
BlMuQ-d�J8�#�E`ډە���h��H0�Ā�q�P%#C��")�	rF4V�}FS���I����PdM�!XA�F�S(j��$ ���N�h;���0u_��o�!�8L;��u�>s���8F����m�
]���y(�	����R��U4(��~��	vj�����i0�<�%�@n>X���QR
��C�vJI\��@�7�s�M�/|�s4n@��恷HA��aMp���F�Ȟ������X���i@B!B �$A��Jl&fC�IPDB�%�\Ӌ��7B��7�	=w�viň��ѷ7|R��$0�M�N􍄜��lȈZ���\-�@��B%��5uCWV-�H��)bDF�2$Ѐ����.��� �%=��i��zV�;��i���$tu{LӔJ`�C�W`����Ce�Ђ��wA��\O�\8����QWe Q{7��0�t��`bm��L�7���>���S���@�"��%W������J��RݡA�E4��mˀ��l��nӕgy�Y0=и*78�\�6 龎�ܹڰ�i ���G��s�F s�twB 0��C��J�� ��$����/i�[��XG�`(��r !+W��NM]Ҭi��<�.�7@�8�h\�v��9@�
π&��9����Uh��]v����袬&;��z�U� �r,Mc�X�hPBT����@��]�p��<*�3iGކ�|#��p��<�]Dkdv`�!�6� �/h���i��H8��{���s�s<�D�	��/-���_k�	�E>9s`�5��!�(ٙ��(��@k>��Ô�.�1mۃWR�s�wѕ�(!�m���7,��ᙄ��wp]����y��m�І���~+K�3ǝ L[yFK �g�e
s���H��}��4u��l���F��1D)'�C#͂fI����|�0]P&C�Lc9��.9�߁�9Ň��t�|/3jB�,�j�s��)��s|�` P`-t!@;C��,K��Zz����� F�(�1ztA�Ǟ�y����ߞ��:���xoCߝ>x�J��<�<�����K� �1��m��8�8:�gO=Lc� ��7��p7�38{3�����ɓ�ΐ.��BL#�&4������&'����~��}��~w�ua�K�t�ƖC�8�|N����='ً~pbZK�� s4\��[���3��"�)&J �Nd�I���  mC��԰8��0Zc���,L�TOG�����2h@�J�3���s/���bY����������~>K�P-��R)ZG�ÍDO�(m��,S԰FkX���o�����A��������QO�_���w/����w�y�U�fL��D���p<���i��8:*'���m�R��ݔ�~�PUԧ��Eb�Q�8�|��T����C��񊚛�Y�h����۽E<��9j��	��;�(�co�i��C�Xmd�	sD��($�˲��
��$z�f\�H�K�pӄSr̤�R��(��6��bȷ6<�a%���L��9F�Rg�(c�T�G
p_�� x���s˄Ж��N�S�j0�8���ֺ���T>���E�;������矃�%Ĭ: ۋ�r-(��2D��(A�z,I棣}��Ə������a�Z4p<�9��c���n��h#@�H�G�8pN�
#��ƕ�ڪxP�@��raa�{�6�A�h`QVy�?�ih��BJ�A�\�fH��4h��),[0A93I4y�r�t�9T�-! �omВH�z\!$����G6!�E z|�wA����-�b@tU��� �/$��;۸�y���oɑ2")	�S$VN:��XA&qq�|���s�d|1����kS�^f& �臁.��@�5�9'�ئ"h �[�rf"�A�^z6�I�x���оa<��E:$�YMF����n��'5h�'�ɉ"�("..�	#O4BCwT�����v"�W�IA��=�U7^�*�\d�Z~>�8RE+���.ބ�	E����^�%�q�I�䂠��N�l�� ,1��=�h��`ۏ*���p��l�)���[B�X�r��&�2Al�a�$F��|���!���2i(��q<>hE���(x��j+AA�����4��aK�@f2����(��/�qQB���1�M>�����)��X;�:P*��9IA�'ý��P�5!+!y�|RD��Bm�VtD�hB¥b"o�w�`�y8.La��g!cC��U(�<�f�. 4&�b�Y���V����@�	
84Q�q�M��Ԛ�qp���#�� qY8����U�"�҂���<J���LsKB���1Iݬ�#��'R@����d�gQ�{�ףC�g��=ĥ:�*�Ej��H�IKVJX��+Z��q��s�nlۙ�[�����_EC�5P�Ӫ?�;k� 2	�V$����w�7���ZκҠl[���9)�`y_}��>'ɏ��W�b�eb�ŋW��T%HPd d��XNc���t���4�-R�ʡ�������>�?G�;
I�bTb-�w^��/����o���y���o��_����=���w�xŞq����+�}����3�x���� r�|ʰ�-t'�4�q���m��TpL�i}�u�#��p��;�K7��MBNPߗ�
L��.O�b8��r!��2����c��!	�Bq�MZ9�d��}����(��G$�<��~�%8��w���'�~G�����^���������A|���}�G�}����π����~�~�_��~_��ӏ����$���B~���5d��e��5=s���������t?�j��_�1	�?��3���������JV�z�Sw�Ӵ������m�`��+pv�cc6���-Jr�/�G曘ľs.�os=�1�(~��_x�׿|��f-�:����$�4�;?E����AΨM�l_����؆�'�_�0������2q�9š[��N����Q;1�i𘬿��H$�S����t�:�%�#:z��]]Jmg_�%���eW5'TJ��TZ{��s���ϗt�q�׋��.�~,U1��6mT��Ȟ#k��|0�  ���|�� ��@ R��p�Szo��z���k�l!� M����g�~��������G�����K�q��o������J>V��t�"K�D��0�IXTcSJ��e.S���,(ѵc6%�=C�����G� ���Oж�斦،�����a�3�n�OJo��}=�Ǫ"�N;B�U�{'��ޠN-� 2����n`FS9W|cڐx�v�h���?3�:=
�Cԫ}7E��8�X�5Z�V����U�jzϭ���w�ޝ�l#�a_5����ta�.$%6e����=���~�.?�5h�Sr�0&�u�]��'�V���n�����F����!�P�RJ
0DԮ �Z�bq(bh��� H1I0L�*D`��$U��$1hN������.�ӹ/[��]K����j��5I��r���L4��W��7@���?7U���`�(;	���<XY�,b�m��V�t ���L�lsLBɮ~�5�?�����c|�*t�Ê1���v�o����}۹���v�(l��J��h�����8�r�&�埂v�1�z���wo+��*|���u�7��\��>���Rj0�A�������|�~S��_2��!}�?����~��}q�]�?��~G��o�x��7�l�����������cP�a�w��/��M\�����s��)��������N�}o�QR���ACW'�������i(��;����i�Jq��y ����O�t;��:��*���=������������o�����8w ��=�3��ZG��;��W�I� ����Z�1��t�\_D����9/eֽnϴ<��ЏPdsPj(���%5st2�'O�)93��y_``���?��u���`��`�FO�"���r����c�r������3݄4%�"|��������d�p+?��/���j���Ͻ��-����>6����;ޓɇ�v y�!�?&Z�t�|g���~�l@#`/��{.��=��_ǧH�ESFȾ��l�w�P3��f<7H��C���x�<A�PTE(��������$�#"�bF�DEPH �KB���++mX���km��T  �R4�T0�4%P	DIED�(ēPPTQKPAKD����g�t�7%r�v�-���q]D�.��F�*��׸����x¥0�qz�E伽��TE��ݢ�/]��xHH�UZ��I?�DL
=��]�%5N�Ѫ��
�P��Q��P�b����,qZg�t˵�h��L"�Pi�gZ"�B�y��z���r��|訊�����F�,-}�Y�H�u��\��b�%��Ր�Qb���Z�ep�]�zz!?s>���>�(+* �TQ*P�kAkA���Z��h���6�(�e��j6ƫK��$!,	ѐ<R2�dhе(���YTEQ��j��V[R��؉[ڌQ`%F����T�+F�UB�-�D�ڵo� �±L����
�ҵX*Kl*#RVUa|�őED0��ʉkF���ZU���UE��֊6�� ����4�"�V[FVڭ��J�-���k
��`������b�j�,EZ�l��5�Ɏ�'b��5E���3�g7~������_�FJ*����9��X������(�N-I�ɵ-�Tf�Qk]�2\��kEL��c�\ ��E�_\k�[kT(�&�`kQҡJѺ]+�صk���S��njrr[hִF+��j�������(�:kAe��cHI?f����)kJ"���L�-��q�Y� ��"*a�h"*���Q�eN	�(����SV*1�1�	rTr g��=EM&��Y�h�Z��T�J֔mi�(�cx�[���+M��G��V����+
���?9O<'�0�Ǩd�c��,}b�%�/�^�^�}!�O�y��Ng$�"�dD�T�'��ψa>[S��KM����֑�$�co&X0`���s�)p�ӧ�S��8X���þW���Tt?�z� ����Ml��>��G�G���@�x�n�^�ރ�cjd�v���}��e`Rf�b �� #61�������a�u�
3�@ͳ�蜗bZ�S=}&�#��5J~lޤ���!􇏉?4�����2<���X&� �FR��}:�����<����薴�98 ԝp�5���l���mC $��fb����#-�@d�, ��w0� ��s߾�n�s1x�p�@Q�N{� ��4��H`׈ �x�@�ΐ�g@�f����������y(�t�]<��؋�����IF ��.�Hs c�ʘ�}Oz����t:�5ϝ�#�~I.%�e��I����-!��犌���,'P����}���D�il��������<��2������1�z8�{\ph���:~L����l���=y���*���/|��E��%>��� �XZB��߇��zN7�{Ï�gG�xp@��B�0���;�ǵ���~>}
'�d���G��c2��'�f8��w���(�D�)@!<�"(����rg�P� �-c��c�C������-��vx��͝2�j���H k!{'H����H@d:��@����l��L,qiG}ϙ��^�/���-��+�8��2~4
��������R��ai�g���b2Ϸ�y"�L�٢�1�ѳ)j�MnM��J�-]z�i��˞��u�g3r]�3�B��"�R�̈P�I�e�C�&?O�(�ߦ�������a�_-a%���{Pc7�לR�����dd`��5Ecg,����$� ���!����'�7�d�Q0a��#"��3�q�ٞ�m���}��G�W���$�����ߏ�RƖ�h5DicK(�ƵmbRE��9���9��9����mM�x�A;\�5&������uN6����*�e͇>��L��
��"�*���N���)��@�6�i�F�ll-�Tx+�r���l��q�%��+�	��k�"�5��&BD���N9�I1D<?���x��ե�+b��9��V!�-"m�u�%e���n�A�)��joo��YSICD�AEIC5UCCCIM5E1m��^��e���y�� ���s��ݰ��-�2x�_��+�Fc���t3�7�yWWN��+12\�Tq ���B
yO�ғ�;W)r��J����B�F��������X���AZ�r�H�"��b�~Q5F�<'��^�e����?YsQ���� ������d.� @ܗ����o�>Fb�����zJm)�$sm����܃�_l�.{��l[VS���ɚ���4�(��-��ͣ���3�4��b�q>(��L��
��C#צ�F�����=��C@ h�%@S'H�����y,���~(!�N|X�@4�\�ҍkR��6"V~`~�����4�/��c�C���9�at�F�K�� aU�{LJʓ����V:_��I6���Y��<:Ҩ�/MQ���S�K(F�����&.ҕ+��|7װ3?pi�=����F�����z�����w���$'{R�����%�(�ru_�����2�v{Ǫ�3"�d��	�7k�l�̅)B�[%~�����S�����WJ�:����DBx����h/�8u*�#��T��E�ۿsw�:Q���;Q�JG�:X p
^'��/�s�^��S�J��Gߍ�!D�u����K��ˤ1��0=����ÃB��a�?ĎK�tYk-R��||�U|o�T�]W�o�#�/�E��i��UU�ב(���'^y/v*%�.d����T0<�[�E�~ߊڥ�=K�5R��t���0�_�i�~]���fa:����|��w��!�PA�"d	�?�RxuϹR}���c'տ��A�f�mR��n?
���8������;�X��a�����y������O��{���y�'
�������]��y����ԏ���#�ݟ���+����ߟ����ܼ��K�|������~�	$ς���S�@�`A�D:?Q��/͎��y����z��z����ю���S����/Y�ͭ����ow�F��������6h�}�>;_�����$ȟ�E�Ix~�NZl�)���)��>)�h��	���v��{VI����HŒW��Xr�p��~���^S����>7�7��׍��]��[ͧ���'�����=����g���_��ߑ�SA�m��t~�������=�s��s�2eUBy"?6V�Yu��~��|8�iv��}�_�a��r�4sG�t}O�U�����_�n��H�H�e����l��O�{.H6�v �O}�U���h�'��3�~k	4���.Y�u����I�C��=t[��Y{F�1� Яd�g�4 ��Rz�O�A�<�i��i��A�v|w��5���j���à��X�� )	O�xr&-��}?F�rz��` /�\#�D��a�>��j3�}Z�}�9������ǧ�xuO����ͅ���ՠJ��)hD��"�&
��Ԓ�У $*�	׀ �|Li�b#���(��)(��彮2���(�.��[K���
�Ŋ*������	S\Ӎ&"�˝n�sqϊ��_4��p�dv 0 YU���(�
K�z���z�Z�Hy�"��~��Tv^x�0�����b�
i���(����%�JvR.�5C�'}��ĺ��Fxuv���ř�0z�����d|Q�0�R�s�҇H�-.y՚���4�R3M`�m���Tlآ�iFԿ� y���]^
^s�W&C1]z9	���)��Jw}�.�i]����#�C��J,*R(ѣ�`_�-}�ཷ���]q�\s���/(�E���f��|%I~	)S�ھ���Ϯ�/�?��.��~���|���'�)/�(������5y���ե!ܽIN�]�h��O'{؉.>+S@j��_)��b�")� �O
^�W��:��싮�=� &�|�[��O���&�bj�:��j�*
"j�����I���b`��b�J(��������C �Wp�p3^8y d�!���q��Ld��D���m��	��Do:�z~z�^�z�� ��I`
jw+&h�<�_��*�/�d�ݫk��^��zO=���h�N��QlK[a>i鍍���j�����Os��:��\}��"�.���V�$�zQ���R�."qĢ�3���h�L
4�9���5�9TS#-��nM��?a�Kѭ��O�#���?��*:�I�̏��/K��0����Gq�~z��E�_7/G�|N���$�<?9GE�i_:�7ףxn�f�4/?�l��M����=��?6N��+��ڨy~f��E|/4�Y�����U;Q�^J�Wt)w=g�^�����~���Y=�c��x��s�����GJpzS ����~�4���Q���+��@�%��������·]c�_C��I��«�\Z>R��3�W��͑�c���	��(nU����oPl�������eb���fb��`TU-i
~�H�UXT��
��iZ�X���
�T�A���B�m�h�E+*�X,�"�Ae��jE�E�")"�FV�ZVֵR���"�"�DdEB"*����* �R�_\27�PRP�T$�13R��QJW^�j�:z���ͫ�&Ȕ���ʡ���0I�ٮ~���d���AA�EDD%��>�Qϝ&x���������������<��}�}���1���kx�!��߃�߿�������ڔi̙�+4&�F%Nl��u���a�Ɛ��9�׶eT5H'�Q?�9�bҧmB��$&>?Э�v���p����~M�Z��W>������ߋߧ_���K�K��U+�D����}~u���'����d��O�C��7��^R�������oG�W��>����D���eM������o��"�p�f���>�����{%�7�K˨G�ώo|���>��x���_�����7�+�H����|��\������<|��ۯ�ϻ9�;���2�R^o{۹Z�S��Uw�W%��E�U�_���Mוd����O2�����қ|�,� d>��k�=�%�v=�<]�+�O>�ٻ�8�s�[��(f9
- �4���-���6�Gt��$�5B�<.�߮�w+A��'Q�w�~�H�xAC�y<(���
��8a���!�O��5��ڻ��T�~Zu���)��|��Rau՗\ r�_?3W�q�I���k�'�P�|r���=�-J��ūۄ��~�^����~�y�p�{��Q�x��_O
"�4�g�S��=ג<.�;��<a�{k����	V��B�X�����EpL�Sև��� ��("``
i,Sid�G|)s�)�*���sP4 �Ǯ�h��p�wo�����+�؆��(t�a�B]�-�Zx�V�����;;���;��ܨ󵤛�Q��)UNvyO�Jw˴)v~[��Iv�ىw��īT�N"� ��oL��c?5�yCԥS���g"q�P��tdOX7j5�n��7a5Zd��&�h�*L.��?G�^ϼ��;2�=����<���������gPB������v�:�~����]����!?dI�a�����}���\�w'�e�29�M%gg�.�u��v��nl	�B��`�Ż�c"�*���ȼ)uq��ڗN�y����^ה*xUp�z|X���Z9���ؗ�ל��Q�v���=ʽ��;[w�m6T��;��
��ۯ4���w~�|C��y�^H�o���l�w��ٺ�����˫�����޾iJ콩ѫ�T4*���c��*ϦF�K��d����Q�'�/����6�O�<>#.�GTE����*SږW=S�/��ʮ�Ƹ�o��,;�x�]�.�����6R/����(8��Nx2���Ƒ~Jϗ?�qپK�;��ߣ҈�N�t��Ӯ>}�A���W!�Ҹ�I{��G���޲S&W��y�9>c�����^�dh�`��.[V��6I �JR�H����w�;�34�������Q�Os26{�>�U�]�.�-����a���/�L��}R䮈ANt��%�7�zl�J�S8���!��7_F�}�7��]a�O���#��r �(R�n��!=����ax�a���Ϙ&,�����)C���~vFr���S%AN��0�L��&�q�O��X��~_�Q����0 �ά&e�����{$9���ủ�c;_�����9�?m���S�ퟏ<�o����p��?����w�Wn�>��ß������5��`�ݣ�2(� ����ሢŃ$�����3�wG`9��UU~�h_�>�
y� 5%�w!�xS�Q�7�{X7��y�b�,��(���GXJ#	���^�I�x��"��
3}���9|Tg�5�I��a�Z�h��G�+���Ӈ�l���A�I���>���� ��O��ګ�(m*|kvM'�?�P�/�a8���x�k�d<O�æ�#�=�'����{(��S[�d��O���ވ�Q��/�`~C�����9�7D\���Q���=nnS�8���xZ:��,9��6g}2a��/�5ǈ�#�8S�a�}���=4�����B|R2��9A(�H�ޯו~p�sg���.����Tٯ��*���>�J�R%#�p�V=�������}���?��o��o���wU%{���]g�����.�o����� �;i����?<�ć��+����@��O����w�Oc�?Q��~��������M@�?/���W0�80|����y��`3�)�	�	��g��z�?Wo�&�\?�Xu��V����??������]	W���0�ve��$.Aؓ�#ߝAV4B�*Х���d�?�����2�F�xp���ahZ�W���/a翇u�=��ѣ��w���W������7���CxoC(>;��3����=�c���_��+���#ߡ�5(��[Ϗ�H��L?�6D����	�.�Ϧ�?b3���8��O�\B��,@T_��?�u�;����f4��1礒���?�lf�}vAG�S�Q�h
,JC�Ky���K����q��ϰԹ/���F�b� s��P����VJ�,*�1�ˀ���Ȋ�4t�j\�A5n�K�|�W�{ؐ5\:r�$�(P�,q�ϸ�oɸ����= ����;�(�i�ƙ�v���C2]�
f���\J��Y"ҹ��4<���i��5��l���NI4��B�i�K��� �=e&3��5�|�LS�a�Q֑��b��"��.��M�J��^d�VFf�IM���.!�H�D�`�NW�����A�^��?�=�������Y�������G���>O���=����axM{�����_���D%�J�
��q�D��>�R��W}/É��:X?�9�CMF�������x��?�Ҏ����&{�6�n�NQ	�X���3M�5���?��FִZ��ŚI1P!U�/�o)��B���U��[]�I󾣮���v��YX�*�U�J,%�}q�lS
rgzUT@.6FN(U��5�k�j�bw ���A���v�.&F�<�
��o�HL6-�a�|�W�Fq���g.#':��`�YZ�7����^���qQ�����I0�x�`�ܘ�Jw���״��r��?�ӧ/��5���ym���TaL��� p5P��,#���k�n��e�o�~��FƯ[�5m�;�G���'��W��*.�*@?RH��i}D~���wĪ�hz�=z�=ݛ/��W�c�-{��<�/(~�_��}f��/㣒���$_��?��eԕ+���=�N�Mؙ�$-엔�Վ{n�<F�v&�O%�Z:�,���%êj��:�zcXj�qIW��-���@� 	 �c !sU)}?�8:����t6߃�䲙�Z"PJ�p�
d~D�}ȥ�����o� w|��T9�*w8��Q��F�y�;����H�B�N$H>�O���c�����A�.���A���uW�e\�#��N���A僔��YN����95�[�\,g5[#��ѥ��6���\��)�����?w��Ɖ��S�=�6f-��p?�=�&;`�����]K+KZZahv@w�2E���:����~���|����������?����&���_��,�p�A�	$�N�hA����y�����/	q�����[�Q���|�}�Z���R��wyБ����/��}���?��4_�q�]��sU�:�������{����������.������k)	!"B���FFF����m��"'��ݫ7�>e�Z�-j"()�r��~'�����w
��3[n�O۹D��wW��Z�X�j�ZXbő��O��}F�elmM�1�6uN��{ޗlY�Ѳmd�N"E�I���qRʍ�kD�����z= 	� Ih�m�ز�RI#�0.	�M)en"�*I��_?<n{ӽ������>��X@J����4��7�jdL<2#J$��Y/�V�!j�S������+G,Չa�Cc!UZ&Zte�cI��6YBBP�I�����щ�4F�F�}]ɱ����#�e+�K�kl���B+����h�,ij�[�{��w�#�dRpR�-J�S�X��O�d�;�B�/����5
Z�l��!ٛhhj��w������k)�|�U������x�7j�y�r���dD��^6-k�v4���b�����l�H<���Ie����s[S{J�|�n9r8���َ���[tA}�v��ޢ�r�i�Y�"�S6Odګm�1�S� kD�k@�\Ӷ֝�Y��>�w������ކ���矎w��w���
��g=�s��ͼw� ߚy'�{>9.݊��6�$��cna*g�|���%���	R:"k�ç�:�~���2�������ag��\s>K�mʣ��_��W�=7����8���W�~����往��k���=���	���DD�����f�cs�������m��~�k��%��PH{��K�6�	D�M�4�\J�(P�e�U])��<��~���>���x�;��^������M˖zvi��k8/���ȧ��;zA�ON�z�y��(͖���ӹ�9?8����>��>c���kϳ�랫��}|��|��B����|3�� ���Z��{���֎�������a�*�e��h���
�����j��	��*���H�����ib�ѩ���V� F�:�#@kZ�{��������?.��w����_ü�z�e����)]VZp��f��)C�o&H�x�0�h��,�!�ؘ�V%��0��N����PSK�� �t��HC
`�˞"Wd�UW��0��6��D���1R�M�Ĭ� S�BRj�qk0��Y�$�d�a���X\�8N&]X�_���Ց"֐Q��'�Io.Ѥ������<ᤪh�))i4N,;_	���  �����c�g�LS])A!.��P�6`%�!az��ˀi��Ĵ�A�@$�|�q�:��:��a������^D9H����eYalBJ
2��N�%Y@��iB��%b"4Q@U��\�'���-׈���J{���l&6�* �j33�TRƂ4"(̙��9wNUT&�o4h�d礁��MU��i��b�`.s�J�H�p�PgH6��)D
28f*��.�h�f�kQ>�d�jѸ��
Ī�Ji���e����Ú5>4��Gh��8@""A]���y=�G��������k�vH�"�)��T3H����g�	\�;ND�<�JXF�$��Ic��Qm��jK\4��-H&yB�b�N��T����a�@�_A.�z��]h�� �^���a��J�3iY܈�
�RQ)�)$�:b�@2�T嚭DEފE��nH��±+��5J���ði4��4�|b�p�ST�F8�I*j��P�)�#���+oԠ.��Hx�e�a-F�r��P�@�G*�b�;">%)��QIWhKX�H�3PU8�bV��~�����Q�jb��[፞s�����/G��Ɂ�S���Yq{��D0K`Ϡ�T@��ք�2YbI��0Fx�����A�tƖ�t`��A�cH����uC��9���7�D�3�Z4M�MK@�=w��QH��P�ٕ-(%��5D��v��'#���J�aa�J��o�gld�`�����E�ʖ�f��^L�#�,
��}*n�1�\��J�meU���M��U2����������"��/!l��/���=2L�+�ʬ
VQcN����@�AR���ֿc	(�bD�Qm��O:J�B!_��S��b*<�P;Sq��y�T4�`�Z�40�*��l^;̳��q<-����/^�zȈ�)��$�Z�-,�V50�H2�	���;{���ck�Ѻ�e�8����ˌ�/�Sn�-��ѹd�kX[r���TI>�͒����nX�����U�`16����$���3��9'�����V�0D-�1-��l4^���:wP��'d�E!��G2˂I�bia�g�cg�M4���-A0�.5�-a��V(0�	N,E����8�N(��QC|�$����9h<ƌq�ZA�/��c��Z1Nt��.i�[HNV�<�3��|F>�PؙS%�/z��}�Эώɓ-ɰ����(�,_3H��MV��(�O���`v8V���0����K �)��2��'���ɢ�LN'k�9`�*v�Xi6$]�_A��c�� bP�H�5�f�)ң��Iy�� � @   ��BJ�������'E�ԑ�2$�`�5Q�쨩P'�<f�&����.��zyɂj"U�����SDQcP�W?q�.���L�A��Bd��#U�	`N��11c������4fQ�of�M����P~y����~��Z���X|��92L�>��!n��`��!�¯v,��#�����a�T�)Ut��b�E��tю�aE�y�̴Nw�a0�ȶL2ؚF�r$�)ffa"����5b2���2H��[N��Y��H�E�nFj(�Z3��v��q�+-�#d�6�6 �ӏ&�j�|	��AVa��vp��X�o+j��fU	�ι��|��Λ�7����vq�a��ˡ�9�='ϋ+�?�w�U��	ϟ*νc9q�����J*�lY��<��3�'^�x	�J>t?��/�q�� i�1���3�r{~[y���7f�+q��-�N�1����a��Js���sPiʋk!+�h��
����[n�P��!B'��e�kr�t�s��D:4ƜAkn���t����{uT����@��'me����%2\�Yi�$��v��D�+�f&գ}A�4W������dgc&v4A�����JD�	�C9�2����1��\n��6����&�T6��59e2�٤x��wDytŏ	'833,)�i0�r�ߒH��,�:ژ��G5N�$>\�W3MF�	b{=oh�ʝ��V������^%/�5�n�)��f��p�	��P�0^��V�d%��#uL��=�e��H,����8�+�}'��\���j���f�S� J��+ě�a=�Q0��K�|�!�cF�ga�Mt��(�R���)FLG��K�v.��j�lYq��z$ ��{=�GZ�U�3�'�?}�J�zx����� �T��GT�ʪ�J6�-��&��M�WS.�6b�ڜ�ڜ���u��2ą
!AKTP��&�cd���hٕ��`�F%� �X@��@M�9��[K�]j��%f�ڐ�u���c�s&&d�ڔd!�C �EX��e[&�1�5+��г`��%Ժ�WZm"u�GYJ�"�ԡ��]e6J:��֪m���mT[*�)sH��[@橵[)\ԛ(�����B�搶J���JsQ[*s):K*�e.�V�Ȗ�Nb�ԋd�a��H�W0.d66UUm*6U�(�9%̥ȧ4���eI�Vȭ�M�l�Jڠ�9T�&�-�l#j��m!�V�[�- �S@�(P RP%)[%���[R[d�W75M�6�[)��i6m�m���jN`9�sb6Uf@��5Q�ҕlmR6UH9��ء�6��+jmPl�ㆵ�ٱl�&��M��6�ض�l%�V��j6�6Scce&�����m6�mQ�+i6D�ʣjU\�-�l��RV�JsJIC��e%�@ڕKj��9�9�����M��[T�-�-��Rڒ����Y�`lKiU6��F��5\�Q̨6
sJLiD���W5
�)6������撮a.u��W5s@lM��Q� �(歒���6+m�sUlq�6��6�\Թ����h�jVI��32 �E��[Ta`����P
U�J�J�"���()ر�EBԂ̒�C
H,R(�P�R�`����i�!hZJ
Z �����HBd��U�"��(�eh�(�
"�ih����8�����)E�J���������`�fV((,
���X�V�B���JZk)\T�b0�MU4�QET�@UCM-*P��14�"R�%
���
q��;����9�~Ŗ��я��7�����?����z�������_������W������w�o��������;�^���u���i�����9���|���z��O��.���g9�<_��_���oO����6N���-E	AM4M@P�R�T��T�QMT�RL�%PRP�2T�-&��0m,V��cb�(��i )
Z�
`��
P�b�(�a�f�3��� �e6���S0҄̚���e�RA��!���)R��**X�J�)�
��X����$mJ6�i�Sd�bf�ce��V�UmM��m(�6,�ě%�&��&a�Cm�M��!�(�6I[(m���V��V�&ȶ�hKh��6@���lR[@�Rl�6R��M�VҖ�-���l؋a-�M�Sd
�Q+iC`�aL�ڤ6���J6�Rٰ6��PQl	M�Y���d�(Fel*کI�&�M�M���U�6*l��J�U)�*�i+i�H�U&ԑ�l�mU[$mڕTٰ ډ���ڶj6��PPD�TH�*H	AT�S�4�D�P�LQR��Lf���MU-���l�lH�M��-��F�6�[l���6�ڦ�l�����dl��Ch6��M�d�6�h�M�l-�6E����m@�&�M�[
ڍ�l-���ԛ*����dX��VS�/���wC#$C%��P���vߋ�����o6>����Ϝ�>g�������?��=/m�>�]W�����/���?!����?���׺��|~�=^?��w�������|�����oǿ��x}�u����+�_������w�7�����W��8�|_��C�&������շ�������w>?�q]s���3����8�����~���^G�������wC�EY	~��d�Q(�v�����Ʋ��Y�S&1��Z��R*���f���������H�J(����bb��"�
����*��"&	�&(�����*"j�"(&)�`*f�
`�bf���*�B
����������*��*���(��� ���B���`����"f�����*�)jb��"
"�
"�"��������)������� �&�������b&��`�
i��J"�bi���`�(�����H�((��&J"���i)�����
"!������"��(**�"""�j
�$���������(�"*$�b"�*
����������i������*"������������Y��`���������"j�$���"�`)�((
"b���j��*
�� �$��������((�j**(���(��j�`��h"�b"`��(�(�B����*��%�"b*�(��"���(�"���������(�""
��I�������"��%�	(()��*"&�&*����*�)�d�����*�*jf�(�)&�b���*�&���j*	��"�(�b&������j	�*�(�����*(���������)Q @H���o����1&����}��8����]��������އ7��W���y����y.o������S�����'��o��xns�{ ��K�!`J �����'m�x�[����~���w������}o�A����M����?��!�/{�z���?W�ձ��_��c�s���|/���ϑ�4}�'�;_x�������oK��o�����N�w�_������B��wX���C�©���,�����r���������1�%���j��>t�y*���VOQ*H �?��E��`�P�q�U'(�b��/	je�1�>ZF��[�qed�������
b�'�L��,i�ӯ:g���9�P�ǜ��I�_�'_1M1�l���m�zU�.����e�-94:Q�L�[D��7�՚�rGE:�\����f�n2��+�����e{�_��f)%���cwf�RJ�2-Q���
}�p�"<��ٺ�����	+FThҥ�$�*`}�^-�9�y�o��S\/=��M��5���=X�\눸��#݃2f��#Q��� MN��&�fX�6-7fϮ$a+@�XZ��&7vhO{c����v�B�����[�i�Y8L+o�:�������pK�iw(3��Q�E�sd���
��ϳu�|�{�&i��M�r:�wݳZ�˴��*����0�T���-���{w�A ��Q���(v�����j��>�&P�'��e#}�)��*L�^��А�?������<��ϵ��L>?-���t��$�@��V�Y��ۙ��>%B(N�R�XE�N~�(O0������MRӄL�&$ׇT��$�>�ف���C�>�C&@޵	9�ed�aP��$�	2n�<�������]���<�ff�a�$�
@3s�œ�3��ό>��S֐��$�Ng5'���*d�gҰ��!*}�}�}�)>�W�C$]�j�������% �2��ѐ��b+^@vhHTGNߪU��J]h(� �J%�@��������U戫�ME�TZ��
��\�Fʊ:�AWYB��\�ڒ�e"�G5wd�v�YR��iM���sUCj�'�Q!�T'Z*W��T<w�U���*�)CT!��ʆ���Qvd-@2�(v'9]P���WjE����i�u�w���9�ʞY�
ʕ��ȰX��`$Ṗ�<�P��I?ɟ�|O���|d���@�BBN��I�|d��:�R��:!�Q�A�h�r���\H��qR���JCvβk���S�Is�--�#����h�T-,�I���d�Me����������������������������������������}�������=�^�;��n�Is�6d�

��P���A=��  <��!�+|��   � ��  �           �    #`                 c��  L    a@����ph&�5[ij�e�EZ`@          �im�	y�D��u�`�h�{�w,`   	��Y�p  ��ITR�z1@�P��b��h�h2��m�      �u�f�    �  �8��4   � �À     ����| �    ����׾   }�    T�����<    
x��                                            	��Q"���    |�8     ��wKf����               ���               
  $ 
� E  ����0 �EaP�P@	�/%kVԢ�����-h��A*<��N�$U� k�O}��L�D(*�'��I��$>�p$T��UHVm <
�� 
:%I@>hv|9 t� �o�(@R  (   � @  �E�F��&�JR��PPA	�     D  o{`(`�����       �0 hѣL�M�$Ɖ�@4hL�=��S��jy<�m2�OLLM�ɩ��m �2L�����&�516	44i�#�H=M�b3S�= ��j@   ё�  �@�h  z�'�*P���P��2m �i zM#OF�4ɦF�A��#&�C�4�`@�2d0��C&�h14`LL�4 �MJ�����OPP�=A� hP �       � 4 �� h     �"h ���2i��� 44�S�yL�cSi�	�I��jcH�50)�`&i����0&� �Mbj%DB ?�
�i���)�FQ��MOiO(�	���m#�P��L��2z��<��4ji�=A��j6���=M��z�Sj�4�3���x���6��S�}�����{�b�!{6��ڮ�R~�y�<n��~������&����>v9E.+���z�:�f:�Gݳ��~�����-�߭�>�>�jS��ra�v=޴8{�v�S�d�=�����Ͻ�����u��������o����'�w�|���ׯ�C3�M�Ǻ��	���|Y��'b�a�w^��-�������z����#��~�x�����g�޳��������1"#D�m�\����q��Еd�Ba�����S�v��W����O��ĵ�l��ÆZg�l�cC��l�0Q�m��9��Qz�U߹�E%�y|\[������������O]��G�R�$��BDS�Mi�H�5��y���-*8s�8Q^�u�Rzj 5�s�����sf�Yg;��4�ȚZva�sF�:g]�����H����{M�v�m�-�b$a���࠰�t�H�2Z�Q0�D(i�z+ߢ�Q���� � ��AT���^=���O*oڟ�,C}0%d�a��.%*����u����U�T�*.���oB�Ҟ	ۅ��Q��-��>'����f��k��bq��|���r=�����ǭ2���(����m�̱�� ����A�4 ��Q�|�햒��W���I��k�"�K2\�<�(R4]����`�Im�*�ND��EO���o�_�1���k�߹����O�(�]�C�{Q2O��3����z��M�/��`>�%5U������9� ��hsTt�����������{�'��zC�z\�� �� E�#�!/wW���*#(�DF�nH@$HD
.ɪ�V#�44�]Ez��Q�s"J0�h�e�9��r�4��h�*ȕ	]�
{ga���հ�n&�(�0��o�W��u���`G��xx{��X�����������FX|�8g*@���������?}���G1�	�x�u�.�v~d��ɥ��R�fP �f��t��rf~nk^���,��EDs1	2)S�TXVv�]z��qAɸ�B��& �`8a�  tH����D'��Iw��gwS����=oC{9�=on��OZ�K�d���x���9�e�l͵*<�@r>縷7h�$��r��@�H��JD3���ϯo���+I�9� 8��#>�"�`�:N��ǀ�x$�� U���X�``a� ��!%L�`�0N�7�c�y�_/k�K�T���T���2�#0RK�
��,X��Oo�=�u�nB���F�!뜍;P�8rٻ]�L�mF���/�N�
�P��ye���I	@C��dYD4`�����x(� ���B`�p�B$�b�l�W�B��l���=;�]	m;�b!:^*�-�H��N��K�Į$@���JZ0�	0��v�Ԓ�?]�����! ���x9�ړ���+�nw��/n����"�$$�d���	Йo�]5�T�g	�vR=x��U���V���U����`(�H2|�b(J��B���b�%�$&b'�@�����B.��@�Ш���L��Dk��nk��_؜~���Y�*3����ɒ~hbt�X�;��"�ɽn�����5pkmM�|�!�3���[E��" `�N��d�#%2�f(E/љك�<@b@P�ڃTR�U?�w� �ǵ�ՙA�1x�E��󉴴�bѥ������{}���o���� DBB���߶u0�
��4��<q�V�(�8�"B(!!�����],$��1f)+I�'T�#)+X�|�R6J2�Y	�35  -��E���L�111� @��>3�?
k����b�٪Z��ŭ����B�����+�� �0I�f&7�6�NwaQk�� ��C�_�}�q�h��~��i]YH/��`�C�VoL_�˂U 9*�&Sc�K���R.�YhH �Jh�5��Z�.�5�a�0F��0O�r ֛d��F�H�DS�Z���3\ �j*�C���1�\���,
L��"���hC0yd�00�% �Bu��}�)�0r�U ��X.�w���K��h1С�l�0�� m�W"{
h9�4�	H[}�u�JB5��.� �$�u\�X�b�ȑD �D��MV��e캚wQBh���#�#�j f�'Pf"�5�[��}����+��$q��N��F��aH��^�j>���2�7�'�X<Z�F-��"��\b�*�bD�Nn2&@�A����@،�:��y��n��U�9ꂚ$!����ZK��pUΑ�b߻Z;(���!��RY�����n����G���<=��G�YiW�K~��ꭝ�ҋ��4B���#;�ĸ�hY�Q�ȣ��'�~&2.�Lc�1\f�r�$��2���0�拱�8�MȦ��w1R���fU�d� FF
��UQ�GR���qs?7�Ѭ �MFĕdzD�d���~�ti����7	�+D�P2bemL\ڬ���T��닌����P��<�G�T�5�m����6��a ~����A��ZwQUY&ـ�VJG�H�#���\��b4�\�s�]�R�dH�ϐ7�'Xj�<�@��xg\��SH�����T|� p�E9JX =P��'�Lșl����K�[�HҚ��aegB� �

���{
�I��B����\R��p��g�2/T.lB�v3���I��m���6��'�$��xdB
�\���+3~�qZ�����2g�=Q�Į�}�YH]g���ng?(o�<�`��@���2��T�@=j�c��*��Ҭ�qd���P��M��������
b���58/"��5�s錡�+�~K��I��!���놌����fC�"H���}��+k��>�o���]\P`o�6�0E��@p�8������n�{QE���V���3p�@�����p�plɢ?IR�6���<�\�U~��?����z2v����\P�U��`Vf��W�G��Ѽ*pm��]"��y��T@ά�{��#A��ɤk*��H�j��f�y�Q�)3z��TE��%(�7��5���ʈ0��UY����J)Y*F�I�]ærŏ��в�Yti�s��UoD�&&��_`7P�6��T}ş��U����,|b��Z��7�RXj�Ϲ��m��Q����'LKx�=����������˵��[-�e0gh��@�����i9����M��fL�"$gԶf�H6$��6Qf�
���O�j����G����'��o?�p A�]�/��&9�}�r��a��Ȝ%� @J(�Ѐ�}�C#��y�[��1�������  �m�R72Ύ����d�`H*N��C��D�J�3����?�=�!޺����F���"E������iȦ/g_|���
�ey�g�o� �K3"�@/-@�S��!�:�w�!a�^�����C�WO�Q� -�}���� !	]y{�!�z�=<��ԒBU�`�0ac��YlJ��Bؐ+!-�?�~�=�;
���("+�N�e�1YYW6x��{�6���ڇ~�~G�� ����/�[�2�@I�M��@��B%&fI*(�<����]xsfX��u#� {�����|��d�h�Ž�|?����\�O�y0��{�~�\��vP��"'�7��Pwm$�[�N��Mz�L�&��u~/��M�C��	�o����s~����g�W�����@
(�O���{���?����iX?�1E��Q)�D����D�ѩ!���P�-" �f6�����MW~?;���?8p����D��?C�������?��q��)uO���Q�F?��&�Fh��Kǁ�!'0��� �8	 �8)��7�9X�D�HD�Oճf��py�X*:<�X��!7���Ѱ"*4E� yF�DyN4�� ܁c�=�F3ផ��X̙�re�j���K�MJ�(��~�ϩ�F���~~��c���ύִN��8��?{�>1Q\y�=>��r~O�G�
�9�TT`��D�:�`�|�&��#%z%g ��6� �d^@g`,���J�+�#	�x�w��	��C����9\�q��g4��q�7Z�߄;��p=)�, c�Q=%+ؓ��i�@Ȫ5����%���Oh����zu�Yb�T�߀�p=Q��� ��\0�YhĘ^p���E�0<��Q��� @�Q�Vu`���W��������ip��~�ڧaҺ�5*��-�����??�HI ��I#�]��z���yR�*����ˀ|f����mxl�q�s>�J�#�������5�Ơ�e礘u�TИ��b�#Us"*��&DO���`Èp�4	�\�9*j
���*�%M�1 �:�$��V�UPwn��i+��J�v�w�t%gmk3�qF�&��wIꅵSLS`Ų�f���C`@p�f�R���b���tqn���cBjn�R�w�*$)�t!RK���팓���E��I�P{����z̪�
�_���Hp��یSB�b�2�>h�f�\��r*���Yf��( �C��.���x"` ��U9T�2���
�`��2������E�h�zB�*MD쉜��O��7T��U˂������XmV*Ve��U��0�X��˖"��u��߯����V,���*[�fˏ�f7^U�
ˌ�07��/p�_�����? �Q�W#�k�%/S}Rb`$jׯe\�c�1E�3�Z��a��v���	Ta�U�,J`g>��8wW(��/(�y�"��b�x&�l�61*��qE���3�6v4�6�(�asB���억b` ��pf�4Cn�g���5wus5MT�Ǔ���E��T��ȳ�=�9�Z-@ @ˉ��ޣP�a���J$���F%,�sH9�*&��7f�ERV�v-E1K�mDm%�}����U��l�̴[#L�|���1��VFgL2�TRL��N�)bRj����������E�Cm��6��l���5����KHRP�{�"���NYEJDP�@D�K1�5MYzm�SS�ѢP�)cO/k�\�@N cPPБL,CMDQK<� ��j=����_w�����_��5�!421BP�R�S����Sk�j=��t�5��ccm��i�)�F�٨S�A������b�ʱC�5-�ԭKJ��5.���wul�L��h�6u��ݣK�����"f(��P������b�Ę�y�5�ژ�i�,�g�+a�ܵP�(���j�(�bj"�D��u�!E-l����H/s�ϴe?�SŻ[�.|��� 	 2������i��[k�������v)��dSn6�yTp��5I�Ĵ�Jd0Z�+RȄa�aaX{�l�y�ti��PP	��*z?1����=�b�m�G��y�������{㻿� �L �O���xE��L����^\1�!�G��H���w�>'�|Z�����֪����=4�km���U�H���#�'u�K�{>���{��w��ۿ���?5���_����������Q���Θ_g���_��佗~��b����O����~d����?�|_\��q�O�^��+������B_�u�L���؟�{�����}A�z�ɽ�?����os����^��������wZ��?��🷲���/��&���w��,��:�5�=��_���?G��'���k�7��C�~?����y�����c��~�P�����_a��M��>gk���	��}f[��Y�wݼV�i��Q�E�X<���v��r�>�h9�)��g������ ����>��nOe������a�}|�no�����W2�߆_�����^Q�~��w����m��W�_G�g��-�V�������茟�X߆=f�_��=n?U����{ͷ������_c�H��L���]����{f5D���?ס�=Ǵ��|�.u����|��Z��_2߉�E2_?������}�y�?��,_������������x~�{"��⇿���2�K�Ogʟ��������s��Rr��@�;��)<Ԣs�#��<O��>9�g��S����8oL���i*c"������S���J��W,�d�_��_�����N܇\�3�1��*���k?�]�!V|%����)B ��u�Z���p�@� X^ؽ����9���q��ex�1���?��_����(@}�|�P��=4������ %#oE'�X{�Q�n��	��U�B����VքQ��Fo��^3L�2 ;�	�B��������ePB��5�?��#���3����" m��V��s�������%�X!|���炭���!B 7����}�}�s��^��q���Ϧ;:�<�<���>�� 	}W��a�����:�壧��K���=^��̿6�_�9���?��?ͻ,�\�����! r;]s᫆���,e��X�����º�B� @	��!�����>�)پ���������� ��>W������}��=  �4��^���|q)Nx���׾�#�xB��?o���ئr�̿���������7�s�E�S]WF����+��/�v��� ���ZŮ�����;M���(�='�x�j��,�f�� �vϷ��  *3������	�������W�>=���=R���c�>�)��9S�=��9���|>:��iɔq�@N�=�{�=�H� }� � @B �����}ǿҋ�1�����ݿ�q�������P��� @�ݟ���*�Ƃ�����k�۫`cK�a���O�̄<�<B�>&�=��<A{��S�i���4�-u�4�(ƲKNG����D�  j��+H~s�]gu�=�������|��@B��@@�o]"��m<��]�U�B��K.ߏ� �/O��[��?�z@��e��m�;W�&�+�@@�*��������Bzv j�~-�?���!$�/�o�?]~�Ѽw��ÿB����;|�d�B�lg��WG���0 MnQH#����<[�˹����wy� ox ! 1��^���宜�����x���A�
|]�QN� ! C��tr��7Ո2\�D,G^p���P�b�_ y�)R��VA��NӅ���|�+/�n��� �ҵ�߀! 4�{ ��{||O����m�����ϼ�X������?�WJ[�  @?Ͼ����%����_Ϭ��۞/����y7��I�d��B� �o�����?!��!�a8�/�ZЄ!�����=����ZQ?H�5@x���l<���BJS��*{o���B���$'�k���n^�����Ny����� (B �@L~Jμ�F4{[�p���'�h�/�w�(�K�V?IR?4��m@@@}�{N:�C�{�W��)�1���{~_>�j�R����B  ϭEW������z�ï�����+���P1Fx�Y����p'�������:�4���h �+l��x�AZ�������K� �0��|���h>&�I�ie��H}�m�� ! +^�4�����kQ/E%���{���F���~m&�Zr�Ϳ>��y 
k����?����C����Y�%i�]������G�������������~�����_J��z���{v�ߍ�mh<��� � 4�8b#�߯��^��)�[�{����'{���/C�ǳ�
z0�����w�w���s�џʱ����RN�t�L|D0J�H4A1���� !��7���gч���q����_,����qa�$-a���?
�����D �P�����L7���b 3�q���ޞ���5H��jW>V�s�6�B}�pQĀ�@�"(1"�a�HHB5I'/bn�E&�*6u��������������ͧ1?>QQ*�U��Al�w��q��/��Kl'�����B� B ��0v�4������_O�6����e���f'����! �?o��M���j�����=����m�.������=�! AT�?���7N�z�x;m�{�����a�tG�ˢ/%	Q@�H L���BB�S�IK�y< ��c��r������*N}}�G�V��_�P����}x̎$+�_�?/��A4տYqj�B���#���ϟ�<�?����I��ͬ���!� @F39P�O���r����?K{|}:��ܹ��L�Y� LSi���'�P��O(�o˿n:�#�ҋi������M*_��#�<}~��h���G�Q�Zg���� ���ǩ�EW�����/�>n��{�Z7��i�� ������_��['����O������޿�h@@�x꣥.�Ž����Շk&~�~��E�-q*"}�?���v�!���Cz鸏�|y�iB,�N��0�#�UN�d2_��ٹ�Q�����bRꉹtu:�Q�ں�M%ke#}���� ������S�!QԱv��I�B!C$
Orj��f]�ځ6�/��}�?��$��9@������ ���{�;�(k��_���R���Y��V����i�������K�>u����'XՍ���♮���|��d�m��%<s�S�������'��_�y�������>�7�Jc>UG�7����Ƨ_nS�8yM~�Ӵ! m��}�D�}�I����G�V)R�4Q+W�?�?�������MI�  Ј6�H���t�Ղ#,�]O�m�:��ȩ�C~�~_O�    �����e�����2�Ѧ�6H��a T%����0��EWmԺ�[V
V"��?�����)��u�g��m�_�.���W|��|n�y�9+Z?_nf|��|x���U0���/z{}����ݻ��F,���*��/ǽps6����n����'���<���^��Ķ��xs\�V��T�����s�U��p����M]��*�������ok�o�^�2�?Y�>o0��z螀�םTg��ߠNuC����LZJ����/�wZg��ڵw�<6z���̡X�z{nX�LP�ݏZe����B����h�����i��Է�S7�ѬMk������c�8�*�*1��{�J��ݘ��e-�n�k�h���l��]�T�jT-���j�R��s��<˼a�֖�OS&y���s�ƕ�a�_ V*���[C�5���~�NC�s���[��ݹ��z�u����v�r#V�z�)�ws�ג�]{-��t��z�[���-�g5;+y���ŭ�h��QaU�Oi3���]S�=֭6�_=�2Q�/z��֧�g"z����ھsԽ̺[K.�D����ȥ���r�*l�a�+s���kʛ��*���.�Rչ���h�f�TO&�=��ɪP^J�jz�m��`scn��}u��<՜�[Q}}�Kٺ�V�!��)�7V8m�Q��M���}�L&����oZ�����
��Ne}�㕚�k���[�u�{���p�g�C�y��K��}V�QJR����ڰ�^�j���k=yt=��-o�����Qinu}��UQ�D�iL��f϶p,;����PiO��U���J��}v�]R�CS���z�Z<���ѧ��Թ�a۩���m��l"!����2���:א���j�չٽ|:/0TN-5�kjZg�ǋ�r�ˁ}�ۊ��zcV�z����2Wl��]y({j�Q���We�Nl]h�׽m��sS���>����i�|��/^��w@�ܽo��u�]��j/[R�����0��}�{8���J,[e__u�������Jכ݌���0�l�[������ڜ�ǚfn�^�0��{�όw�8��wj��W��g���lú�V����gKSԬ��:��9�x-���={jy���=x���)֢�ޭ�؛^�{�&�ړ�e����/l��m���l�J��cu�,���g{�	7u=�+�o�N+o֩���u];X�Z����r��7����͋n�{��zѴ�zvkV��u�j�ڽ÷�:sGQ`��^L1<ʎ�a�=��L��y+��Xƹ��+��SW������ǽ�1�޵���T������OZ�oe"ʷ�M��{{�"f�[��[��ֺ��u����:�sj��;��{�yeں�s�b����u�v\;�+G�Es�gn�WSa����ǹ>�Z)W���j���ڊ��Su�i�
�iY-=���ws�uϓ��ʝ��u�s��/5���O_w:�
x�cu_97u�
�v�딸v��SQ�g��&lն�}�tPN;qym[2�W﬜�F�Q�emh�iN�7��آ{������粦�/��^op'���>]CZ���Ԣ"�4�b��L�v9�mB��^��b��Zj1vq���/���۸���ƶw{�<�z�A��wS���(y�]rQe�Z�)�/;%׹�N�l&i�r�,2lce.��ط.��j��}��Uo{��:����=��]v�O6�m;��2�)���[Z�Q�{<>gki�W-�z�{v�/=�;[�7�	Y�6'��5�1���~!<�E���G�k�����]g7~	$�̞��|HC��V_���:�����־$�ݟ>7˳�co� ~�$1�V�-�����R��_�� C�"�a
ګm�l���:ti��~4�j�e���UDi}e_=�u-ۘ��㸳��Ub�ci�G�b��g���䛛ݷ���j>}��L�E|���s}K�Ҝ�T��wqv�J��]�nh�*g�,��a�w:6�5+Ke�����\��0.�k���p��B�Oj��DuF�]|���t���S�rv�]��Xy<�R�7zӳ8��xqR�]�k{���j>�ܙE����EK�eTQ�';�}�dOj{���G��EE|YX��{��a�s�y�R֪um�ە+u���{viW�5S�Q�F�sv��g-\�.r������s�<짽xT�*�ő��3)˜w^m����E�[_�N��V#mm���iU֌֏^�>����}�/���w����J��:�K{�nT�,���˭�HS�c��k�J�B����]�*:��{���n6�3V�ڕ��.���;����*�myާ���S�ek�s�io��<�%5�~���B��Z��L�\s�y3�ZlSU��W)iS&J]�/�}�kw���ԧ�S��Z|�W�y�ﶬ�7�^kǩ�VҘ�o���f	֣�ʙL�Z���0.�#���_h�b�KZu�R�*[F��m{vW���r�u�+�ml�j�"[V7ɏ�9Ȉ(T�o�1�Z����љ~/���wW��'����Y�=�Ʋ�x��r��)��[�}�S}C"J����>�ʉ�¦�VM�0�ea��E�V1SK-FYJ��)b-F�Fi�8$5%��-4��#(��,aO������Zv�i�W�v��KQj�~���){dN�1�ܧ�;����r���{�5��4=�nW�楴�;�w�2��:ٹR�s��{wy��{�\[Ne�s���`�G�/�L2�벋�S���Ԧ���_!���`Q��W#��^�=��<�<�R�S�f˻�u)wi�k;�ϏxO'&���U��\�>|�Tfj���CD�}k������5�ו7�R�7��z�A�/�v^���#��\e+|=�[K�*6���5�z��ި��j���Z��Z�j
fm�c��MO]��;�.��>�����<��{�K�b��ǵ���k��]vD�.��/9�S[o�}Jg�[�R��G�ي53����Z��ʕ"��K�n�9_�:�*�@��r_u���=s�Q�׽|o=�ᝪ����]��w��u-�k��)}�׏k���d�g�,�gP�bv�qj��iR���V�J؍j�f�Y�vՋ�=�^GZR��k
{m^�En
]c��:uS��׏{�/���u/Wk5��S�E'�����U�2y;ݔU���x����²���9��G֭j�ʗ�8�s븫�s܊�����SjV�j<[M����"x���[4�|�MTMk�{��շgdR��g=���*Z7m1�c��np��u���޻������h��Nz���s*�>�&mma�mU=ԩ�u��KJԭKj5�h�|�{Ƕ�U)�ƮJz�=�G��z�عK�u�^o"��a��{7ޕ�Ը[�`��4���3ח;c[�ps`���\���"53qY��F�غ��^�v��.��iF�\%�S��׷����uɪ^�neFd��+[�4���=�w1F�n6��^����S�'vks]h��u�X֖�.]B��3D��m)�i�{u[�_{ٴ��%�Ŷ�F�ufiG��Z���w[�^N�S��2�.5m�*��{�wW��wz�1�S���z�o�f�&n���G�)���v(���2��٭kF�T6UcmV����i{nb�m����֮L�%�S�(ږ�-DE}�z��D��P�o��iŪ���S����j�h]Z4�Z[h��Vճ&���أ7��zq~d�z�&�֢����\"���Iy��֢�{��/��J�F�ֺ�%��./�&i�c���K�94J!F�;mD�4�+{`ػ�p\���5es�7,���[n�l�KkjQ��c����b���)�O<��if��ԥN5��{l��E��/��{�*�gj*6��A��m�)���D��Um�*Q6����V#���^�*|߽�>����Uʢ��ZiF�YQ�Qjl(��ٚ�|��ST)l�eҞ���mm��i�z�����yP�N�έ��0�E�Ʉ����ڙDPPT��n��<��3�[Խ�d��>�3�ڧm۵Ҧ/޽�6_J��'�]��ƥam��u��)�-�^G�oS>}޾k���W"���'j(�����Q�9�/iu���[f���׭֧b�'�U�|m�����}����(�o5%����fּ:�L̪)Z�Sk(��덚ɐz�R&-b�ݗr^��m�i�ͺ�e�ۺ�k�ZQ���Q���;[��#j�J�:�[,���^�^+��2�.6�k���f<й��m�>�h�������<[kUm+iR����]��y��ɔb!m���)�j�<�ѱ(�Ay�+��.�#-�R����}j���7�+��MK��"��kl�JZ\R�+|읃!��&�l��-���Jv͵ϭ��BƵg�9n��CF���J4bV��u�a3Km�&p�*�Է��9+iAMq���h�D��3+:�L�Je2�DIz�Y��_qU�m���p��g��
�)y�=rrQxV���qSl�x����/���k�9Z��j/��mU����KF��\ާqg9<���%��<Wjږ[m|�U=�E�}�g�ڪ����Dա�Q�c�S�&%f��6��vئg�{Z�/�h�[�O6=ݥ{���6U��)�͉D�.�ǲ�sOZ���B�2y�*ִ[kD���{Y��bd񮱥elj��ܞ�2˸�u���o%Kż��֡���<���-ML�ڷ��T�U�v;��S������u�u(v����./��:ѼS��%Oۚ)ו���J:5+k}�uo9�FТqih��L�,-m�Zĭ"�۝�������2dG�ޱ��O:�L�]Kϙ�K`�[E�vΣl�����Mo>��g3�^�[��D�`�ټ�W%��{zV����jz��mm�Z������C	b�����
�SS �31�\�'`����i���5Km֎�j����._qNPZ�j�kEY컞�oR��S��b��57�#�cp��n�-�E�57v-�=5�U��{�|����:�v9��ڈ��1j&J�=_Y�6��/��N�U�N��v��a_vu���v��ֺ�{�.�DGަ�[{W"���uٕ�PX��y״;�j1^��]K-���V麚&�݊W%m��R��vh�2���o�f�k@Y�ku�7[F��L��5�ӝ���ќֵ�[ǜr(�k�c����,/���(}J�U�B�oԻ��Z�޳y�sso���5��ƥ����ԥv��oz���ރ�Mw��d����yh?@��l�w��[��)Q0dmRW�a8�G�8-�L�H ����_/���_S��ݣ��N��粽�o�����r�gc��=����������������*IpQ�B��HT_ﾧv�k�=s��-����m׈�d}�O���[������Ib�0��S}x�6a�~�KP>K����T$XI�f�]H'���m-�_��wsn7������q$8��R��&�.4t�q��8��%�z���\����
�Yi��1�lT��3��gO�L"2!bմ����<d��fu_;��X���!SO�q�S�e)��șb���\�g�=>\�A� =�\I�xL��"I�8%AH�I�)�N)���cE�r44�i�rT�����O�6)�k���B���b�E��қ�]>�V(W	Lv�@�Dp$K���.�~�0�^S`�pĭ�V��T�&��2|�kr700����秽Bk5�e-,�eYt8
u	���.4�:�*��ѲF���X6�}YjB�QYR�i�\��v�2�=�zl�47#�_	h�c�UB5J,qH�P���DS�_��40�Z�ut��;�|�4q9��R�V2�7$C�qg{N����H����2�*�Ÿ�&c+]�&��S�{Cj�������4�F`z5��ZT�0���|�G��V]�x�&��|�ZS��Y�j�c�i�R��'ŏwP� �n�Z�)]z�b@��#W7Aؽ�Jecؿu09��?3삸��>Eq�Q-UÐ�w���4����I�=Ree_4����T7�����K)�d�s��ͅg�nInr��
g9�2`ۧ[HG�5^]�a�V��5TM�Z�f5�V���%�=�j�s�xu�ei�0>�L��HZ�A9	D	u��5q��5ZY�Cތ�x%>ɝ���	�����|D���	 JW|�p̓��ͨx����:gQ
ס��<����HE�x��ͫ24�Rm����V+D��[�6���*�4�1�X�D
��	�W
��`G����IȺp)�'`C�M��U�-��Y�*P;EX@�J΋f��1�������3Ć�B���cW�XN��b�����Q�ØQ:�n�)x��9$�f@�C:ˎ6��NiNj!d%�R=V��AT��fp��k��m��Xs]7���kl$����CJX+��p��9�(M8ۉr�gV�J@�|�����7J��N�n�-�e]���/w��ݭ]�S�@TS������Cۘ@R��CTD@�UUA���4Q0�TPU4��4D�Q�MP�L�PQLT�T�QJ�"D��UD�HQ!%4SI0DST�JPSKQD���GAi�:%j�6�7NPIV(TS��Up�%*�TW :FK
�Q&�s?��2���@�O�{5��0������>��LO�����3����~�M-8����^��y~W�?��A������~����go�����}�}������`��B*_�'��ϡ$��:��21�`j�V)�Qf�����0���ל��|���s����l��gO���/� Ե5��5tPX�r��U�$o��`�c� ��v#�I	#�Ȁ��s�� ��ƪ�"%W��)��x:C`6�~"��I]1��5����hv��=��K�����N�\1��{��$�'8��4�/m�2+��@f�0w�e�'	�������p6�A=�M�,i�ƴ�m�xW6V���
�yXT9� c��%5;��%w-��G�9�)�4�N� �ځ;561!+A�7���r��l���ˆH�]~�()��YvC�I�ys6���j<u�%oZ\�l���\û��J���OW¢)f�($��'&�O���@�
<�F��V�X���KǐR9�$�!D{$�@�3��ō ItT\sA�l�¡��G���*�A.��,=J.�s�A�6P̿�������'� ZK�@ܸ�~��(���1c���x��T=h8�~i��k	dNk�{qia�t��Wn�2ulD�-�C�Z �X��B0�ɤN?��/U:w�"&F�]CtU�I�|��C�]�Y�l�Gv�;�ˁ��r�J喍!A��`�8���$��n	�`��s`:[ɇP�gm[�Jv�b��ƈ�M;'fq��g���,�v�0�C��O��	�R��kv�1t)d�Ƃ�-�e6�Tqs���@�(�y4�X$Q"�9�5Ir|�����	���p�����sR��k�,��3yL��h�o�2K4��`ع�`�k����v1�X���D�DQ`j��j-�UZ�`e%d�Ί������Dr�4ܧ��[s��U�<c�D�//GEO�N4�c�{S==8y-��-q��%��i�H����P7`R���.�^ݾS���dꋷy�x����E2#�:18_��,�TG�5y�i-_�� ?.���b��_ln�['QzM�q�5��ڲ��+ =\E��C!��uB�1�]�;�l6�-?"��]\��aT��<�:�d��a8�H�*m4��M�7��y7�Ӂ�x��7�Q)�Z��q����,@5�J����j6$ea���=8�{������nW�����0�x�8R��bFW)9�C�RcTD�-�{���ų(��pvY ���!3�Xy���$P u���3�5��o�%㬈��^h?=��(O�q	C��[5S	m�i�=�(I=Xq!@��K ̀�L���"�4������慣H��
��*mr���o ��kj�^X\���N��c�*O@2a�B�����EZ_aJ_��O}����õ��A-1�ό�Z-��LLz$�
�R�c~�q���@�{<1D�}Z�#���3
zͭ�6c�;�@�j�pQ_���U{͠:�����׭�x{�ʄ���e ����+�T��a�`&�$R(/G��y~?K��=��G�����q!6PM-A��t�T �����P��Nbp�4*�Ob!H�ƿ,�����~_��C<�A���f�Ҕįx�������JS��(@�.�
���C��b6iM��h{#��Ҡ�����{�L��0m!�E<��N{ܙ��������m�-�@���`60x��ԃB�JJ�Po?SW�?w�{=�غ�u+���1��3y�+�>�mv�Q�oyd��&�6`3�4<� *"�h��j���"����*a�
J"�(ih�V��j�b�
ZH����*���������*aJ����.}�u��=��v<g�޴m�Ɨ��1���v��h�q��M�ⷽ#=���GO�&��[������r������,��K��m����������)�O�����Ą_���@� A�Y��O]�]��v:��ŭ��)�uv������k��W����������Y7�z�:���L�������Ư��8��j�" ,>���!D!�����O���vҰ� ���S����������!�,����$h�y������z�g�I��_�0�|x��   ^��bAn�`_ᑂ�G$�q?L#�4Q dR�?j�ɘ�~��F�!�H�e�����3s��M_>����q��1ttOl�%��cZ�˰1CC)��F���p;G+�*�v�?g�π�E%C�N'~es��}���#���}��  ���M�h˼s�޴;�/?��N�V��  � b�J�HЯo�oa��i�_��p[�����Gq������]��]v��h3�EB�%���K��.�00!�� �{*?[S�D������u���o�qu�.np�5��9��,�]4Rtќq�L3-�M�=��MUF�K��Gx���K������eU>W�S�Ӡm62�.�,2R�%k�!�(��ft��hL@�6���/(�~BN<�.�3.�O	����i���ГYs��Brh��Ns�����FgBUq��\W�S���пv�yp���9j;�y�;��q��,�<:�Y+amho*�Z:iswO	��8W�?���_w�,Ԕ�V�B��mL��cm��PO1Ew(�'�Qdvf�Һ.��<��B\(�
K�	�#���d8�y�<��z2zT��G�CW����JK��Ǒx���,zc��P��;�z��Ó����o#���؊fm#fi��3BT[Z�i���s�M�(�L�R�%+�S�)S��(@	Y��l��Fki����iىq�c0�M�V2
@f��P0% ��Q�H����TJ�$��l�-SA2R(�*�!C�)�	�Q��o� He�f�)Lͣ`s�k�����;�l��1�0t�ͳ,J�Q �L��FXJ�h��q�]��͡�Q5��QP��D��-[V�]Ӟ%&���Í-�RTE��� H(�y%F$E��U�)�ň
S���P���3.�W�;�8d���H���	Pc��������&�B��������5q���^�VdXA�?&@QU�!6�<�bl6�N�m�
A@\�� ��R���l�a�ƕ�T�T����98�CCS)T�Ra!S�j"&��I���ƕ�`� ��C*�A���[��q:t�TB��
�Z*R*bAhR�9�(ULI4���P؍���������3��[���G��t� >�@ "�-��sP֜ʓ"����1I�%�9��l���*��
d[JI���|��i���,��R�����H
J��V�mP["�T[[R��x8��P���+	;����^F��npI$P '!	��,'�!/X	���Q[� d�Y["�FNH8ʍ���\gN\RlR�ĄC�C0��:�$�:�K�(�l��$�G<p�`q9H�#�F�1��W)F�����%Gv��E��R�2ڔs���tbVT�`0	��p�TR�<���L��3;�Ǚ<�+*Ys$�)�9-j�|�u��<�ݬs���O0���I��ՙ��羵��omk��M�y�!-s�{��������w��۶��
w���s��/9�u�a\�K9(�+x/����8�������d�B%��Ϸ�~}�j9�T}���]o����>+P��l[K��y:��kLj����.*�}o��2y�u(��~�j��R��׋m�*�-۞S��U;������gY�U׺��"\2��u������32rf �u�-^=j�5/�ֺ��wG-Aj�.fǷ����D�e�|<j�({X�X�	�T>M�im�����g'/�����N�Q:��F""��f�>hc��;�|���v����z�W�U]��}l����(���*6�>b{��Y�����x�z�'%`�Ŭ�{{�掅�R,iV�����L��ب�an�����z�Q�D��\'�y�}v�ȱ��!��2_�u����_��vK~����\���\��}�{�wݡ�֩��k>�_����Q��m�On��ϯSr{U}n�h��6r=G��ϰ�����>ra�}��Ty���.<��Fڞ�)m8�R��_�����7�m�kN|��>�g1c[�S�k�Zy���U�_����q��r:��o>{t�B��5����_��z���%K�#�L�i��b��f����r��y�����8~���{��}�,~=��FӼ�Ck�5���fg#:�\��#��X��ҁ�K�0�>�މ��7�v��uoj<�������_�:���
��ƣ�Ub�}�w�&[�W_���O'k��m���ػ�W��z��ԯWi��X��6^�����qki�a��u�w=��%�F5��As
��֚��f����/={c4�f�LR��R���U���i��N�����hҵb7�N=ze�_�{�o���w���QyS�ڈ*n_p��4֥�U�v��ɐ����b��B��`�}D����|��+~���c5�{�,W�������}N�F���]i�뵿v�b�^j��W��16�޳,sk��R�w���~��s�i�92:��l�7)r\ߚV�V��c����m��wp��+Sb��-)O]�Zu)_o�M��=G����6��x��N2rl}�z�N�����:�ѥb�y�qk7�<�Wm�}��)֫�X��Ԫ�����'b����N����k����'�k�lz�S����4���?7:܍O�񅏭}��f{�k�[|�����ȍDm�q�̷����GvD���m��o8�����ܻ[}gn�L[De��J�y�}|�_y�ݽu�P~��S�����{��4�4���kR�ߩ�=�kײ�(�0ʢZ��]���������/�wL���<�y�5�_�d2E:مi{fw��ޭ-���n�9!�m��L��TC�乊
,�eL'���-g�7�⍍�(����Ä�x�S���zУ
���۷}�1��ڢ3�o%��v�\*�o�}|�|uQ�,u\�3���qU��ֵ3���SU��Rִ��O�O5W��â�l��=��Ŝ5̧��䧪%<�\�ך�S�6��D���k��5.s��K��}�Yz�녍��e(��E�2�u�l}ү׵�u�����Uu��QXRԴ=�s�"}��j)���>�բ*ƾ����c5����E
�[N�Rh��T���L2�z�m�"����wLʯպz�kͶ�u�>�����+6(�;Z�8|��,E^��J����f�>��}�1[S�{�z��u���z��\��M�~�{�۷�z���Ü̫o����V�:���Z¨φ���uv
>J�~F��$L���N���m��q���յ��gjݹ4���^y�[�O<�Ͼ�z���QEb��V�a{�ϸ��gu�ЁRf"�T&d��N&����]��MM�<	D�D&iWD��2%r���C"�RV�HedXg��2�A�W9G:��P�Ժ`y	0� ����~2E�VI��{Ry��r�2y'� s UΔ㷄we�F�vb:�v`����~��b�<���ܴ)D���i������{�s�+c�O��ߜ ����!'�$$��\��KPTq{B⥓5�f��564�F�:�d�d*V,
�X�F�J$�T��$%)�$RP���HI
j*$���(�"�ihLT�1@PHEU@QC]�P�# uܽ��^�c�vc1<1���a��b��=�Փ���f	�uI�_���د�O���:/%��~�"��7��j�f�*�:]���{���ڦ��ݬh����������~ö�N��}��������#������<w��������oI�;/��}؏���8�i���:sGz�?���/���b.�An݆ >�J����m�7�;�������G�����qO��|���O7��o'4�b��L�c%M�li�^G$v܎������7��[��6��ދ�뵃�d7LdQ���k���K?�]���Lz�K0# 	�F(W[T�����)�;m�h�E�fϩ?� ,��y��\����Sy����Lq�z�)�<�m�v}��ֲ�S]�^����� BM�b�A��10��a�4ȯ@H���T�& ���.-��-��T�Sd���d�})V��c?U���$����C���l��y�Q ��q���`�[F"��� LiǦD��6˂�!A�5��$��n1_UЅP�=&e��(��+�%I&�2���G�rIy���.2;��⇧0�i#�n��7��G��[����8�����-�'�6zQp��?����/��t�*�c��-�;N�&%(}i�=�9�b�2$aS
q�	id�E�DX�Ip @9>1w����{����m�
��B��/�$���0~�A�1��TnZٲ�
L�3�$����=�Kj�$mmT6���H[@��q�.4���e��"mEiX`T� �
DFY�q��58ӍT\b\j�b��%C��%��6�
�aQm%%�
ڎ4q�!m(�F��E���M�%O��Ɯ,"A?L�8�F�I �����9���E��{߫�_���("1Q���ZvZژϝ���_�ڛ�機Jj$��fN*45k������X���1�q�qj�hk*e����TՄ�8Z�:~�`�)&@+���1A��
���EH���/3�QgR�irdT[��?t�GHʊFFu�x-r��5Q�y��׃�r�SHR�	���
C���22����D�$HeP����7���J����E�Ԣ1QQA-�1�b�����$��"1���J"1�`��%8�ɴ9�ٗf�l��6�$&�|��u�2.Q)3+X�J����E"�AsSRV!mp�QQ+m���m���Y�3��ۮ�Z��%Iu9&Nk*́%d�		�N�b�y�EX��u�d�(�F@E`�U��ɒ��l�T
!J�5���ADEsEb��Qb3��DE�mB*�F"��QM�@Рb
D	R @�
�d���̕����*�(�rTX^���*�X"�&�6�*��i(�j"*��bKqA��c�1b��x���������g+�~�ß��>��ו�^��~�#�������\����b�I��GK���n������~�~t��g�+7��\��^�9���+�V��g_[%y"��Ym��2(��X�Z6�������Z��`�,�D*Eb�R��0�#)H�Q���! 'g�όeP�PUD�W�޷n3p�t�N��?����Y?�t��\�!~���m�RT��G��,�~��6�e5�:j���|�ȭ*Jo��\v��M �^�?�%��� �N/_���ڝ�4�B�����0�
P���␇�d����L�d��ʓ���)ҡD�A�J�Z1UDDV����T��!mQDE
��@��A���Z�`�5P��0��HM �J�b�k,��`�UU6��Yl��sS�T�J"(���u��*�����UPF(�`�E0��)@9MӁ�y��8�������n]����yN|qY���̔�� YH���i�����k̎9:���u�������:[!,�vbT�0ħ���F�ւ9*�ɭG�/؎gM[Ӹ�C�'�ue=E��@��;�8f���"�=;ώl��&F����Җ��e�׉9�ry�]'�d&��L�_�B�h'�K{L��eg��_O��T���)�i%a	���p�R������8�����;�YZ���2�<�FnU�n8���߭g)�*�}׬u�z�+�W('F��`$���� ����֊kZDZv��7�X�
Dc��B(gk��s�u
s<$��h�l���	��4�\zA\��#���1�:�6��zU�T+%�%#������[
߼i2%��He�Nk�!�-�R����a��{yǰ�r��+p���U��&��,CJ�\߾f)�U�~�s���6�\��#�<��8����춀�,a�\�S�8�S�LX.#w]�Q�UB�M�4� �eu=�����Th��?S�Qv�#p�WI3P��k���~9L�?�88�`����~�(u}�n�ľ0��2��h*XR���,��ne���=�f�� ��5fv��7���ǽv��M ���2Ds�SG�%,�ߡ3ڌ1Rw��lP��E�7f� ��d����B.�L�[STx�_����6
f0u؄�*+7��c�	q��8q7��Ed��H��%�P��������%j�gRkx�ݮ��7��MՌ~*ׂ]��u&�)*ѢDz�
�!�� Ǌ��N����I�+_{�o�@/�+�w%�M���/M<n�ob���s��m�i�I�^G��＂5ҭ�l�o�����H�F�.Ĭ��͐���h�̐��͍*�j:Ԝ,�k.��N�qOj;,�o���4�v���!)���B�g����r�>�b�"Z��C��ͩ�w��T�&��[#���r���bX��u<j��g�;�*pp�\M����`�[����b3T&'j������EA��I*h�h�=��uB�q��i�"`��{�����Ǎ<�p#�D�i���,=��`(����QK�4��ˑ�E�Q��yVdsl0-�D���B&A�����N%���e�A'�ȶ���|Yhј�]
]�"F�h��sE�����������B������pR�	�!a���*`D�)(PX�Gke�?���c���.!ͅg�hE/�/���N��*'�K�X�}k�<��@�9Tq0hU:�dQ�ߢ��A{�����OO����ڽ������ە�x/��z����SUA� 1�8�H҇)/1 �aRÿ�y+��b��V2��F(*����
V��+ej"��
#������U,bԠ�؝�d���Y2fE��d���P!��@䒦d�f x�F`"�>�U@D+*�ְ�"�`��b�gZ�"�b��1H����C��,U�TX
�((dbVAd�m�$	P	�`,<�*]��ª��VV*�Q��eEA�e�*�,TT`,Y#�kb�EB�2/���T[hE��4tԶ:�WfoZ�.���
�>--��-����TQD*���(�,A�+Y:��q�M!�U�V,X/���z�]M��G���`q��,"��;�QR(�UZ�$�&��

)&i�)����"���(3���F�m6��N��s���ZZTX,cl��E�mY�Ff����U`��()IEUc������K��^��y�.o���}�������}f��Qe��~����$0�<��))d�S�����	w?�t@��Ti���t���"����/�����ۦ�hgd�p��Q#�J�ǆ�O5��miL����6s)^#-ha�)�{L&���6C�L�	���1Jć#ҙ)�?��\(� O2��;`�S�8%������	,c�΁���alX�,�%�6��t�9�L�-ӯ�db�CylG7��I���R�Q�ĸ�}����*,{�	RT�YP2��l��7����1ʇ&�q�SubneK�0x	ҧa>1A���	�H�s!Ewmp���Ḏ�-�"5�I(R]^a��S�ʱ�d�3=�aE.FW��ky��EO�c�My�V�t�ϋ��?�����yY�A&�[����q	q��KD׹�r���G�j@�+���& i�4���<\�9ᱏ�s��W��X�D��o7�e��T��U�I�}�*�"���ʎ��S��nخd	Ce�"�4�l#�Vw�8{",_.��Ԣ#blQ.�̓RP`�(�0�k/q�~�H34W`�/%���s�q���*����G�|��<� s�|]M.d	\@V$��X�эK�nJ�e�	��\��]��2��!Q ��<�1���a�?I�QI�-�Ye���)ÅF �6FE��A�R%x	/k^��^�c����N8����l�ȡ��ƹ�*ĪicfidMv���pu��g`/�>,�.��/�&B.g1��y��8���ۮ��%�&nH �[t�$mR؈6�4� �b\��4[�	�� ^鳄�����.�L5"����O&�w�g�ҀS�<�Q?Ȫ&c���P�/3BЂ����C����*Ar�=&��i3 CE�  ���J��]��zחZ���&r���3F	�u'@�S@���Ke*�P�S(O�Ү5T�Cc�P�踸EQF*D�[j��b*R�*5�*ÙPEUC5��`��敔PX����ٙ9S4��. 1"Љ�e�(�jF���"�(�iTb(�*�(�X��H��"�@��f(�Y �*)�%`��8!?�2@Z�U�e֠�d��#H"���%Nh�u��@�kIT��a�B"i*�*��&������EQT�H�/��L��2�ȵ"�)$F�B�2sB��`�%8�M2M-E*J��b��G��d�Ú��f���ybl��(��4cJ�,F(,�b��~_Y�-�,G�>d�$�A`C�6�
�y�2�PF
�ȰEHd�5�#�"V|`)hJSA&3ҌU-��*�)U���Y
''�&O0�������FZi�*R"���1�)R��߇�??3'�*2)
��M�E�aY�3���!��������,�~~�Ox�b�)�JG)�Ґ�RR4e8�[��Yw-#JW[X�eI�&!h�ih͘CZt⌤qq�p撐"hq.�`r�+4�W���]�G�����60��k�[�c1Z�Բ]��c�/�c��L���M)�B[�����������DD�M��F���~os��4�-vg����*������{�Νg>��`C������f�������e��5M�h��F����bT�� 
2 ��'��HTBա9��-�H-2m,�*�
2al�րQ�Q$��b�T*8$CQT�1`���#0R��m�%��X�F�)Z5�kaQ[AFՍKK
0YX#%B�m�[KeY`-IP�%h�ch�E�@�(U��[�*Vm�cR���Z��g�����-)%DjkmX!E�dQ�i[S��(
1�g�ЅJ�$�{w���E���C%E��,���:�L�0�"�H�X�VEDd��
��4&&!(��F���v� ���9�E�"�Z��H�"-*�%b0D�O��H� Ĵ��R�4�����X(�YU�X)�
+ P' rHd��u�h�cHQCKU!@� �� ��Z�b��D�D�J�0DP̕  �|���
����-��*,�Z2*�((B*� �'�'�MW��""�Ab0bJ��G�*̒�XJ�&iDġCAE4�QQ�,R�!Y2���	�s��+	*By<��X()5*0TX-��E#�-%EQdzьC0��3 Y"�$>E\�CY�EP�RU4�H%�iB�a^�V(������
O2�)�+�($R,'�J�$���IUPU�������
���
�a�N2��R����St�-�O1��d�IQZ��C7YE�aR�*h�`��V0�B��.R��\� �g���"�(�1�)������e* �$�!�����+Z�X,"�$̐��OH�����+2V���Fj��֥a��$^J� ��a�92,"�
�
���e.̡٤8�GgU�m]1�-!P����TER
���Y6�L�E�3 �
�dAb$��
�E��e�IQH��Q�_6(!�	��J���l1ƛJl��j�;S�K��lX
AJ��`�$*JȨ������AL�U��Z�(��X���E��Hve�V�.�	�v#�q�j̊�d��^�E�e�
�(��0`�#�aKmjV��$�
!+d%@���!�R,3cYX�%`�������	�I�(�AE�kP֨�R*(+H�Nl��E"�d� |�!� $��1T�AE���V�*�b��+JE"F/�eV$�i���*JbTIZ*��"�C$���[)ۤ�ʲ�f�7,g<M�
�V)�T��1X+l(��*�K`�`��UJ�UQUEb+�P�Y$�!� %@"�T$�$�<�X	F���P�Usr��ř+ �Xf
�ml�j�)V�,-X�������Y8���eiG4��LA�4�I�� x�
<��B�Z�!XJ�Q�6�c+
*ŭDQQ`�bF��Q��
fdXE!�9�
� � B°�T����� �$��eB��a���5l*,"1�ZDF�e��`���A�12"����8�)�s�-��Զ��T�P+:Ձ�+�
0)i٥�+E`,�DY�0���1Z�F����1h��Q[aTb�K���_�5�Z���ɔ8��.��Sb��+�+��`�0�����YB q
``�&�q D-+���RVQ�m+*�D12�R�HTSHM$EFTR���dQ� �%EDA��������2V�-�X�1Y-��R�1��d��((��PEAb G���)H�P���<I�Λ'�~����y�{^o���Ǆ�}�u���^w�<���y>���3�zOY��.�(㸴=��U��o��K�����Yy�_�@	��&�3a��4�Z3���Qv����|��>ߌ��n�7!�o�mM�,އW����}���a�	�k�Y�����~�B}�����o�/�3B�-���DX��CW���+�+�*	�?+�θ?f�?Gs,S��|�)Y��Z?4 |(�7@��9eR��=�4i����΂&��r���卌5ģCT������T�S*�z�~S�E�e0m� y��/��������:�,����>���M�.���`�[Enk�.����q���@H�uK;.C���W�+��G'fڴ��T�/�saq0TR��)�p��Fo,���]�����27j��K4D�f7�ξ����A'C�F���OiB���u�u���48�<�)/A�Z�cPצo��Q�n@��0�3�y|m���ZB�P���Iq�@�^�Y���^��K
���ij��@�u��v5�'NN��L.�R�D{w��y�R���j�e�ws�[x� ���_}X̱��V�b%s<�2k���+�"���Fu	Ʀ."����l���Ү �
$f1�G(*�P����ƕ��|_�Ӊ׵� ��eܨ�GӋ/5b��6<��+�7�Gخ}��oĝ�
���7雎9��w����p�ȕ��g�D¤ESeztCSx�ׯ�
n]�U�3��2*����m�M����!������|y��`�nuT%�q�>��i��*�s���n�l����s��˿u�C�Z�ȕs����>I�-U�|P���S�� O �+K��LG.�)�h�m-:w��8�k���#q��*�B�<b5���h�,8�v���FG�.����I�>��X�v 4Q�T )�������;��C������F�����%���yS�����iQ�0s0�f������dt*��-�\��mV|D���	sҮ����p
�K����B�i���:>�ч(�BrD�v���G&�lY�h��<�TS��s�e;b����9�:�w�U<����t#����l�Y7��x��I�_ziR�
4������h��lÉ2�J�(s����rH�9��iݦ���%�����ĥ8)۲d�/7. rWW��C�cPQoi+M���F��?ABj�������#�K�+dH�T*����t�F�~\]���`p00ک�{�3" ̉Ǟ�����)����� �$�9�m�m@:##h��]sGÅP�e��\+Wr=��s��E��yEe�cS�Pl�!�cp7>�6W�����#\6�;R]^�2ϡ���3�]BR� �bx#�wS�ɹю�)�$ڈ)�`�`T�K7�W��.�Z��mu=#Mk��X����q̈́�g�ߩ�q���J���`���1c]�.�����h���׫�H�K��u0�� �V�`�|�`1}`Ӗc�G�dj;����A�eN�������:�,��ӊ��@t�s�����[Ț�^`���h��<�Z�u��x^6d���nSk��y�����r�����gos�K�X�oN'�������c��������P����,_�}�z�v��'���o����~?�
W�/�	8�T���f�b�o��V�\�@9jxU�� �>���K~/ �� �2\��7�Q���Əx�(AZ��9��Eu10�-c�Q0.��b�;N|�F�0��������d�ߌ _�4b�b(��v�QaƸW�o4HVW$�Pi�yբ4X2F��=��u�	�}".57��v�V��T=*u�l�Q������=3f���nHu�`��N}�N˔8Y��s��H��$��p��!�l"�k6�9���\�� ��VN�]z*��)���Ig�13�uF("�Y��-R��5��wQ�h���Ep�&��/��kMA��9�"	��+A��_�z��!C\��NR�(G�7RA�A�ôXG�a�e%j�H0����9��8�<0���[�薭��Dc(��*#�H��h�c�����'TK��A��mޅzFJ1�Bk�����٨��N�*����I�J�4aڹ3���)l!` :��g-j�8�P���`~��l�C�Q6]�������i!�'{�ȸ��`z-�V�Ҋ2�<r&�-��zck�4ΐ�7m
؉�UE�9��Ja�55��TQ���\V*�U$��*2�C>��#. �`I
�A�UR�vv$�1U�F�&��T[BWM�ә1<�kF��3M�)�:�J���b�9A!O<2�kd9��H��
$b�"i M�@#&�^pF�d�.����)�Cx�-2���z'��f3��$��X�����������_��_��ߨ���������R"o�_������U~��x����B�mw><�dQUQ�CIMI�JR%)BSS#M# 4%-!EAM;��j���t����X�Gm��?f��3�E#1C�)"��! �R�cT��ڢV�1�X�*(�HH&`�)`���E����h�'�F8
�j���C�C[&Vbm�flڙ��)�T�,F� �P�*�X(*�P[a1m���[AI�]�~����������a��)�?��>��t����/���	�ri�����~���W�=7��A=7���&�1�,c>N�_�ôa��Xa��W�E�G��$-���Ʃ-�l��تmm�KeU���j�q�M�=7ȓ�K�����Q�eR�%	E��A�t�kq�:��}��~��F�ϖϾ���?�\��1�?�k����>����#8��r4~�.��o��������w�\�6y  �@����ϖc7�����p�����R����k�� i^���˙�*�3��!���3�4���^��y���q�֤�Y4��W�w�/�(w�����6(b�|�rƞ^^^@�     @���Fth��q��"AZ��iXU2�(� ���oq�@	p6�����&�ߦ�>w>j���~a�4�Ç6VK���oU���d�(��;�� �7�{�
�ϼ��s�_M�o@���eD�-�rs�&�y�1��/�S^�:��i{d��S��B�C�` "Γ���HWI��/ Y��>�)缗���[\�u�&�{Uo��|!�W�?2h��nkM�T���@��گ4���Q6�S2��u��+T�H�*,ӝ�P��k���V!gJ��\-�w��d�װ��[e u��8�3��8��ts��c�ɦ�5����l �+[
d�c\(�rЕݥ���)�&M�|,9n��E{�^��J���η��l�������*��3C����|ñ��o�} �HЊG`�;�zVc�`c����Ƌ�IEN���z*��v�=\���[�v��I�I�2���T15��R��0�=\�?�� ��^�u��s�UD!�Ss���9�p��xH�+����c!�kj��\J%S�b�X�Kѕ<�������"ų����0�%�]��ި�͉�[�ǱPR�X��=R�i�9|��3���EM�G���0y�W�b��*���8���D/t;�L�|<l\Y5ūe�d�A�uf�*���(�-;C>���Vnw��7���i�w��U9�2��u�������7�oA��h��j=b��Ȼ%��Ԃ�����#����h���M��"Vi'�#����r�|�o�y� �����٩r�2n��.iZ�=��~������Z��^Ԩ���ؓ;j���32
VXf(���;,���o{�4u��4���U	��8{��d���i����ŏl)ށ��}��ʉ�E��27?��#R��	���m��̹N+/Iű�U֓�bE�x��{�����.�^��.���1�ͬ�!UeqN��|�$'�"��'\���5�&=�gV�
#�4�v0:m�]�uH>D�0���	��)���n���1Շ�B��(��	Q����a���A]�WŲ2R���T��C:?ήX�iE�.�Y��Zeج=��o���Ҁ�{�tpӓ{t��id�+��Վ!0l4���ђ /l��0�V�Q>0"��K��7��gxk��1b �|-]�X��2��sM4H2�g���Jt]Ed��Ve}�=��Z�OJ��uu"Bk�)��sӼ��c�b��E�u I��n�_�s��=NB~H�'&�-�~	�mH�k���Y� q�骮qP���4c��'��N���b^ :�?�p��|����v7�n9'O��>�)�$J�
yO�7^S��?%��y�.߱����x��l�g�ic�w]=�����?�9?�;�����(�8���/��F�0���ܘ��Ds��5��u���ũ!P������[y�d�b�yB�BA�}G^?��⫎5��ፄ���8`ej
��+�@��t �R�4���,&("G�D)�R$�9O#�m�"���J�X�̰}��N�r�V#�D�:�aV!j)Ȭ6�>'^����hu	�M�➇N���>��ԭ�k:D:�L(�¬�CJ=��%���T�����v�u�:T�"��A���Jd�R��`�v	`[H,qQ��34��K�T��4q����G
�"��C��m�@��Q���a�:����w(����l<�B��>	\��6q`k�*��_1D�y
}��8�2�%q�'"��A!�@�$���e� ��J<�xC�6������*qVc֞r�CLr.�fA�~8�A� �A�l�$�EH@Q��M"�Є��v$�T�,M*ŢAC�aU�fx��S-��.���9�g�a>j�����"�z�V�@��&!.�0T�����9H��q��
��+��DW<*�BI3qĔ��ixS��A�#\�F֊<�V�h&p���9��	cn���l&�P�l�KՓaq9u�FH  �����UpW8�+,Oa�8P��:vDNC&�z
(@T�H斘��4�����@�z�U��,��@d�sj��k�I��j��E�>(E����e�"�a� �	n�\DMA��DQL�� �kʏ���2�����褺j:��!�:W�⒕,��8*�\�h�
�m�IY[j$) ���TTD�+X��V�U���(* �[�QF,/
�4�P�X��EES)$�$L�K@D�)M%%P(A`
,��VTU �+
�"��
�
�@4F
�T(��"��Ȣ"��<��}o�����������x������l~�9�W�ucw���:O���Nӽ��'���/��
uk��l`��^% S�]	 @VU�A�MTD�Q\C$L(deTɊ\��?g�<ߵ����=���~�s��{���i����xP������3�×�|����fo��� B�kg�=e������^^^@�1��~s#������̛��	�xE#2�3��5��8��Ma7_�@�q��$�S�|��n(��1�->`���diVY��W'|��~bn���n1M����l�����*�� h�<GM�����7���'x�(�8�.�Ñ���֛��.w+��5|����y�?M� ��C0�
�x}�#�I�;�G5|n�*�9����Wϒb|�;��~��	4���N�F�T� k]b�H��Ĩ�b�ɞo\��C�l[L)�ȗ9���Q���zLw��8v��ٖ��ݗ���<ĥ����b5bu�c��Oɣe���a�˪�Z��?�ns�H|�;��bl���ΆN�z�o��O���D�u$�9��Zp�N����Bk��y�����{�/ �Ǧ�f���K��u2�z��uVˑ��¸/s52b�R��.�]s/u�]������[2���q�?ZUc滓���O:ȟ�J����y�u�P98�Ql7@�f�R��%it	�bˮR�i �c"��B>;�u"QL���e�>��Fc��%��0�@�2��H��$�6����[��"�1"-��s-̞>KJh���t��On:�0��W$Ҟ�#ݻ�݇��H�9��x!���k��f*R�G�,}Ǥ��O��xM�S��OT��4l� V�K����]�.UM���`W񏋑_����8�q�BN���
�e�"���1�ntŝo�Q�02�o�H����)k�</�r�/\bC�WQ�Y;S�x�aucX��D�cF���O~2�F��a������j�I�?�)���+�����g��E,i�ge��{G:2-���uf&��|��东�Y{R�c�䱉k"�P�Tq��Cޮ�q�,1�D�yx8L�Ъ�a��"Y=�)���Zc>t�`U-��L��H�]^V��z�'� �O(��[#�*H�����r������1O��PDs�ȧa��0�U�x����-b�y�A�:d�hk��d�E�W�f��(]�(ƍ!d�|��FlcĬ�Єy�/{;�ǎ�����k�C[2^��i�@Õ��˺�.�q�.4�e�'�C�"���[�D_$���㶋1)J�8$bp�.q;2��G�'����{$S�l6��X��@�l�Ewv?bvE�Wb�5��g�6�7�ו�t^O��J��1 ����ȧ4$�A̤J�Pޘ�<_�{a1M�&��y�G��}���f7���^����F-������ƌځFd�P�(]h��jFR'��BH���%�tY�|�f�v�x��p�J�~�#��z�s,� x� |��x�(Ϗ�h�@w)r����!�_F�%�ku�����Cze|� �  ����Ay A#�S
�0Ż����^W�z^���?G�q��g��B��|o���O�`��'�O�" ?s���{�z���g��|􉑕�K�i"|Ϙw����v�� V>a�)�Ӫ��B��T���R()A��o��"�8�D��@P |�F@���Q�cjVD��=۰�}�)"�	@.���*"�w!$�-Y��aC�g`�Lt��6�d��ED�M���<]A҅��D�*�Aˬ x�`۰$]�ЗU����7�2ɒ)�Ib��5w�ϠD��5�Ũg[��`~D�PtUE�S�%A�tҟ����xs^AрI�^�H��̨�TN�փE�@����"��`1��l��];�
�W�+���X�QGtP.N�LR�h�eA��diP����X��d�6�""B��ɪ�8���փB�M�`���3��-�yJڢ֐֋hF�3GE���.+`�A��5b��)�D
�B�sŨ8Ӹ���4�DR����}N z�,5�Eƙ�H����8td���3BqΠ�c��{F]Z�������M�i��r�B���]e1�A�9��-$$�U�	3H�����3K)�-�4Ś��}H^��+S&N��$�D*�J�4<C,�4 v���
��*�B@"�H�E#,�#왲lm	]��R�!�F,3N ��`��p��(��霭謍h��D��TQGR����y~tr���Q���G��}u���?Z1��RVF�,-+ZTb�Ȃ-*�*"�c �4�>;��F�SfcfC$�E�U�E�$�PX*��(�()�))fJJ"JJB�� ((C""a�"�
}���9����7y�=�s�_�콇��+W�x��=�_�|�t�^#��M��꽇��~o������O2y��J�\�K y��߁�>�s����E�~��$����ߓ�?��b���%#����sR��I�"ڹ�F���Q�񾟜����� � ���b�(��������8��IGz_%.n}2p�B5a	J��g���F�[(��c�O撙����Z:\��?���3I���n��է�s�����4�{��$�j-�  <�1\	�����U�ԵzC����Q'�*P�D��M�_FX�6L�1�è��p.�X��3-�t��W�Ev����v�ի8�i�h>���q��+�]�E�d��2�1!��q��p��y��]��O0?|߅�.�&��Ġ,b+�0g߀���h�����\Xy���	�����K�̐
N������>�����7.��Y<{��~o��|o�Ǚ3�Hb`�܌���m;���ȿ�w�����
C,�:�*o#�w/���UY������HT�f��c=,V�u4K�D����Cue���B!Z�5��ovu��c��7I��ԗq�����6i��:���4t:cuo:������cX����*!	_�FQ��-5��f�U�n%9^��ş����nΆ[�%�_��^w���>���'� M��W$:��8���*�E����Y��99��ֳN�@�����%;Y���{�F�q��Q���^֥�y=������NlG4S��V�ÚI�]r$�'#�����P��o.��F�^�x�`�+�9t��L��%��9�����[^Jy���C0��c����B7l��\���J?�Xz��iB�͘�2�"����S�5Uң]��F$K��D";<6����oVu*S�|�ϔ��J:�óx� ���=tM<����M�\�ꥯ��^:Ŀ;���/�¹�۲�vv����n�X�"�I��'ӡls�ƜO3>f�8��`>��iEҾ"_8�%50��d�s�6, ��j뚬�\�p��~t��gs�L2Z�P7AOvA|@!]Ng����Ѹԋ��z�:)��Ӵ=R���ٞ��$�6s2�!Q�S?���V��� �+:g��A��H%��C��HV⍈��nF��:����TŔ�����a
�/�86�V�:��|���]�o�܎�%��5������	?�N�b���ҽw�}����:U؉I�(h��ћ_0�N_1O�E��}>\�=,Bz�Ik'�&�N"}���<�P�-Z�xwM�ev�z��g5�n!��"H�2���O.L��z\va�oi�1��D�F-(���P�̿0�V�m
���B���d٨瘙�ө.cĔ�}����w�K9�׾�␪I�̰5�	��N�rDF;q��������N��wẞ,T!k��Z�Vf�3���Dk��z_�,�FK�U3!5h�8�['�tPhW��s#K���«1콍\��Q:r�ÞJ��7Nx�}������������FJ�~�C� e`��CU4\�[c���G=ؖ�6M�U���b��iK$�R�,���/ 0y �U�}x�W�O��`���~H���~i_�|?��G��e#�J?1����ߌp����Z�,��w���7�G�ٞX���=�IB�T ��a��8��x���
V��g"l���dfi���8�а@
��744F��E�����$c
D��pQ���
a�Z��ȍ�O̍&�\r*RD��sRyAT�H�H���J�&%}GB�R�ZPͦ�(|�e�z8�r���粱υ8���tC�c�!*�'��k*s��E� TP���$i���G�PI����0@[� c������s�` ֩�R.��EX%��HO]���� M�i�i��"��/xK�X�WP'�%x�IV�N`"Z�WU%��b��
�Q�N�u�x��^��#d�I�LP�u�� D�hP/)�@�j� B����I#��d YlPĎ8��8�/4�,S���h�"(�(�Ђ����` %T]�Y,��>1�1 C����I����Ď���Z���H��L,�i2#Dc�+@��$
��e�e� X�g!YBY�`�bFL���h�$�43h� ��,VL�N-I_�=�Ju^p�	xs&�𿟖��.������1���S�~'��%@��YzB��6��4a�6�[2mZ��c`ư�QK���aU��(q�EBr�(��Uj� 2��,1EHQBR��`P�2[BR0��c1�o���s����3b��XZ�+P

IRҕ$D�()���������nS�鏹�{����ׯ������zG�>ǯ�����ޯi���/���7�{����8/��p{��1���1�*?BO�������+���h�N7�y�5d���5����#լ�����:Ɗ��md��On��eOhOA�=t���O��PB��k9~�6{�ofeV~�gG۝�t�쏥��j�VZ8�����u��y L�踙|�r���2!��n�&�2�m�Qi��|���m��J�X�}u�K�|�g�j�B��f����k"@Fa�'�f��yB0��Y�oGw6��S���P�c�4�$f�g�K��:����U{
���b���=ӧKy��E�8�̅�w�u����J�
�l:��{�n��z��4�|�f���s�`�/� ��Z;[Ұ�qD�#\z�9�[]LL^��j��`��}[�f� !�:UV��D��˅#0�Qq��n��[�����t~=Q���   �^�=����g����������/o����E�H�����|WK�=�����������+�d����?Zg������K�/�o���1<�_���s����O��ӛǬpBg��QB���Zr�R�iw��K�뙨|\h�(�����W*�M��WM�F�{qv�E�A�7>R��>�Ή�W����K0���.X'�@�>�&��6��^^^@��jeWI�abEP���i+�d#ӉGWGU�̸X?�0����x	�6U�[2�A$!Ԯ!��ȭ�1n�}�o/q9�zm���wI�F����߸k��o7Xվ�j>e�\�T�ɋ�������z�i��C-+z�>	
�����-=\�]�5!��G��7�L��S�>�喒���9�r��B�+�ht����BNA�;@O�:�y�]����$�
�%�nXU�Υ_oRnle�Xz�~[62����qV���d�#����6i���Z"D��)�t�����9�F��9)��3�N�:M�Ez���ih�����]	d_e����V�?Q���c9��;�� 6'�,�3��BK��oG'ֻ�y9,���,���)T�t�z��>�8J�Mxr�α;�q�(m��.�;{�ī�>
x���C�AÅ�N�Tn����;c��u�E'��W�}�T<K�AOg������G/�@H�)w�K�t��\o1�_
�BL�r%Q!��b���o.����D����rZ�6��fe�ݐ�3�ޙ��S8�l	��O k�ߛ<T��� s��	�i4�����'p�gz7 �ú�tS(0�ͪ���R�t��ϋ�h!�����!���&�dٻ~FWa�@�Ao�ŴI˻ud���l���.�H/>ƅ�����0��ZI�q�a��[��;�@�L�Ӆ��j/^�Y�VS= ��Т��8�|�A���1r��^)�$݄�u��V����ib�L�-��'�ƥX���Ρ��JI�E��ޘ��t=ef�v/L�g1�Y&ĺ3�՘�yR�O.�(�ܲ�U���C۰��u+ �i=������":��l�u�'ag���.��$w�&Ѹ�X�x�$/�k���Ԧ
�'�g����fR�iNp���S�n�#`ӖB��v	i��r�,�-JK��_�����X�e�K��Ꭶ�"Y�ǹҎ��)%��e�.��<�ǫ��dg[Ms<a����땭�+��8���S�#CFE���s��gJ��+�#�D�ӹP�y1��vjL:8�2�k��`���6�ǚ$���=��Ȱ�5�O�5�3���5�r9�A�C�!!rGg6�i`}��3�Xdv9�����LY��u������"��N�4�&v�@w.g>r/S��
Y<��xr��pZ0���+g��<�-���9"����IWEu5߱hn�˹љ0�`5٢�\&X� 4K�|���k�`{�;�7���z<IZK��ny��o�|D��z<������pM����#֍s��R�%�"C�^�V�A>z��!�V&�����  yy�|O��=x����z?P��������g�%�������j���չ������o���8��'n�������ï������f�\M"�g�&��HM� X��0r�X������I� 
��)�*	��(Ae��b+#����Jq㖢�����A,{
�c�@�	$ (Í1@K�-����Z�2�dB4#�� �163H��FL&0����m� �y1�9�r� ���JE2A��F��Q�����2��y�A
����������g�}���\[_��݉!'-��Z����՘bJ(�PȝE�g#"Dr�
*�i4���`�0��C��$4Y	�UwQ�y�1F!ѝO�x��� ���:C�9㶺��d*����F�ᶩ���1�P��b��Q��,I�xC� �l��	!� �z$��F^��J��N(�,òE1P	)#�*�� �*%>Q��(	> ����.	�����L�QB���в�́� H�"e�$�)h�|
+B�3�@�yA�Q����7�U�	zq�8"G8I#ZY�:$�T��1��`�Ns�H�BY�d�=CD��]�IP(�pa�6���^�ס��ԇ�=���!�{y��OC�u�����Lz��ϝ�Z��rN��g��D�	SyI�XJ�h�&�i�[ZU��1��"�C�(0�I�
E�� �hP�#L��n8['���3Ka��
� +����u���<&�*"�W��?'���W�����������>qR����Mo����iO�U�/ y�����m{
��v���&�O�D0��Ѣz�qx��u�rkXA|���m`ضDfF�I�qs��gE��f�H��k@F��x�qq}�/��hmUs�Gq�����C��h��[��m�ҩ��g��^L�#�q6I��sTX�5���J��T�S!U��Z	���JV�{7����3j[��q`xT�(�⡘�����G.*�Nd�B��'��@p��������w�T:�dg���ID���f�D]��{=vZ��ݮ�=J�p��B��N��S��c(�2 �}Y��;��_�*p����;�U�u5��UI�P�e�Tb�a�����Y�B:��K�]��}[8�'}Ա`�f%r$
!S��BJ����bjŢ�] ����On0�n-��&`lغ�ri�!T�I|�[o��l�*�Џ��~߫0r�T�����ѷ	e}����s��L�	7��/0iW��n�7hؙڮhn��;�ܺ��8j�5�l��06�r�0u^C���|������9�� �N�n8Nl�f�6�*�	�Y9@Vz닧�n���ݭ���F��m��s�r�y���W������ˑY{���>g�O�9��3Vp�ɜ݋fèO��ld�dQ3;����P��e�j����.k��,�&�����p� �H�" k�� �� ����??��>���a���[�>�����r����z?�_]�{�@��=�n}B\�f�f�~��}�=O]��c�	����B�=�,����r��s��7��������&�=(nh�J���^�f|/�+һ�6��H-^�ݪ�!�%H�����mŹ���~�*]��N~�i	$�ؠ<�"�����i;>c���k�Z�� �"́�Ex|��3n����2���ְ�0����%ݎh#}���ԕ\[x��G�Ԯ�%�s���b*�K=�ӼRwl�q.��Q���Է���?3�@��H|���F�'Ce1��<�q��:;YG�[_����{�M{��<X7���ѻ@�����"��
	��Ѐ��X�O��*�iy��k&�3$�������=���M����,��R1�n�Bu:ui¸���8HS}!��d{�arl��.�z4(�X�q�&��:���)��QZe9�E���Qә7WΗ��&�F�R��"	��g|^�?ȣk�L�3����ȥ�k@?N|�+��q��k!�{;�`�|z���z2�8��_�w��5�E;���d��HZbݹԓ��Ӽ�q�^#4;�E����D���O_���9�-�7h���[�?	�/���r��R�R�f��d�eNN���rf�� �/������������D��=�wN�xr�[u;�U�
҆�"�اd��U�"�
+>�N�u)H�^��h�v�7v'�����S�
+�.Z%x�#��H�hb	�#m2���<k�~�(:�����D�!�Ŷetk���sdiWLB���&�0��iUŋ��on���Y�M l�>���r��ӷ6N�ɫ�:d�vD�eϟm�3A(�hL�A�:)s}�t)�_����Lxj"I����?r�<sG{0r}�>_�r�d�b�zn�z	"KiB>u%9�_���-�k�:�oz�y/2z�W<2��b[��!���>:�XJ!I8����J��U��.�F�齒 �-$}�dɁ���o�+�n�эI�ֳ�<	��oLM���x��y�1D��+Lq�d"v����o���B���V�i���e�b���R��5)��Xb�o$_N��?�}<.O	�=�Q���3�b-����J˸u!m��c�+�W�2a	H��>zk04L\�d��'ZW��2},����^�����͊��x�]y���55S��G`�S�9�Wu�0�EZxP����7���Y�����/��=�=�����G��
�.c��������v�pٕM��V�$;�%�����O�|z�b�낡|��:�eQӦA>��캑�}���.�U������f��	�_Ў�
���\:V�
H-��EZ;�]�J���gtZ"��o0�R�vO�V7ì�֔/$'{�m�������>�V���5g`L��&C4��*r;�$��pZ�2�t=!5����K�ۛ$cu�=�Y10�Ӛk�Qq�T(3|9�,��ln�{� څ���P6�d�d��J��Vq̽d6�=�fz��C;�Q����� ����OG�z���_a�|O<_�q?�G�L���D���D3��S�Kk�M���Gj���Q4�-�Qe�Ec��=��������I � i/�J�v�\A��G}#a0���YM��+
��P� �����/^����g'�;����>L�lv�	9W�t����X�Ͻ�U���������I=;���\SO�?�Ǿ��~Q$,���EǙ��%3�R��S��4SB[N!�IW��i���{_����e��x�i�?�K�UX�Ǐ����N�p	��,��mb��Oi"�Q��g�R��9�����~�}s�����}5����0c����v�a>���.��<�����N�Q8`L��H!@`πA�:4�(�)Fe�t(�_��7�]���Ͽ���TAj}3N~���I�T����6�<���o�4 d � �p9a� ��#�!��c�+��d.�LxM5�����Xs�!XQ&�8�c�F��`.8�PXN��O���� É
I�k#,�!�f!����W�x�c^G��!( !�X�
�s`ޱ'��kkm�2�K�kT����XlQ
Dg�����US�f�
hiB�(�2�iK����|���_��u~3���?�ݻo��?���<f��8������_��8���P��� �bA~�8��aq�*�Љ�1STAđU#TS%DPDTM$ED�3UL0Y�H�
Bȫ @(#�p��]���8���\��w�֗=�}��(�g�i�/w�?`8=��{�5�=�N}���l�ڙ�7�^{^p�����%���BrB�������W� � n�?�Kny���l�5�$���tB��j+ְ�.g��%�3ȏ�I3��������j�>�8�B�Uu��Cw�3�|�kK�n�c�f� yf y�  y�yyS�yn�"�Uq]R�4';{�p���G5_�b��	���eWY�-�џ&$؛Ppd�x��̍��$
�D�T��e�|Ey�4ம7͡�CAKz����$�b6*��g�t�O�d� u�.�9&�z܇`�ʼ*��eg@f�Kj��(�P�[ʾ��	���b6эtMI$
��ҿ>P�T���C�� �V���LUkp"p��A^�t_�E�ut@�WH�Z�����/��̴Ar@D	9j�O,}9G�xQ��,_���>��!|K�O �ҕ&�O6��o�O�q���d>�iPM�E���аU��n@�d�Y���%�6,�����@5�I��!��x0�G��V<
<��6歭��<8R�=μd:�_E�6K �aGČ���E��]�v��IAȺ���,���/F	9�Z���j	W9�!��̏Ʃ�6��5�ݠ�|y8qM�V��b%_V�-������~n�h�4;m0��d2�����-���%X"�b��pY!�Vը ��dZ�o�a�BY��A��=nBһ�lV)��X��)�R��^���,0O9�@� R`�C�������v��qyӏZ�#v�,N�5z�h[r� t
T��&v���|��wƶ�ib��} G�;q?QF/
�j!8 �\�`�:oud���6Xq�kFR�_\u����5:��ʡ�/���0epfpO�=D����F�Nt��1�KE{3��]�b(�"�~��IW#�j�琛F��q炦b:�į�h�K/I�&:Ձ�OxIC�� 5��Z�-7H� sw���]f���ǂ�����Ze� ������9j��4Y�:�+����f�;6к臂�?0�GR�����3G�0Q��a��XvË�U�V&ݜw!%B�K��V�X�^��G��"&t㵢[4��&�a(��^u�7Ä�C=v`^\B/���_R̒P゚f[�����L�mǮfPj�]�7�ԉ����8PD�u�ڴ⸲n�]�Ā�l�+̈́���I�e��bi��� �	�#P��Ug^�7��ʩ���fD�<�W���UaA!��Xz�����%ω�7Pd�HC�AP?K�39��0�*we���Q���tƼr�f\��ɐ=<����_bٚ�)9�*�O}����+�I�:v¿G��e�ہZR�2�ּ�)�Qc�si���ةR�a򞵁(�˥��U��QYJ����������%��p�����a.KVhMG��8��M�����"0������}�2�WHA�C��[��'��tqۦ�������{R$
@"H�����t����y��0�fy>xc���i�����W��w�� �U�כ�Ÿ �x�0�4t9AE5��3�Ğ5(����g�4�>:��o�]��V�y3<�Y{�Զ��<G�K���=���7O�oh�o�'w>��	�)��:g@��ÕA5������^*Ϧ�9{�����t��o^%�{�Ǒ2�8��>���]�ƃ��-�Ƙo��§��ߤ�_[c�ի��>}o�}�)�ֿ�d��Gc~r�����C���K����w�٩�g�_o?�$>8w�%>����͵>L�h�q������Ϝ�b��M7�}sD���	%�^1������瘜�~���W��E}�մ�E���o�6�W��=�{��_Y��f�x���/x�qۿ������H�"b����������M����>mH���?��k���_���on�8���ǯ�1�"�. �5�f�1K1E.�8��2%Z��@ŉ
�%B�N
��1�s�/��=W_���c.C����?+��������]��u8.�v�?o��|��9o����+�����hܻG/���?6Y�h�q\V�[O,h�<iF�����[X���am�"�k�r�Lޭ'����Y:�P�Y�-�}UH��n�B��-2�~�<P����q�_��gl�]�Vn�u!��b჊��hΞʝ9
�S�lC�V��mo�WE�۾��<غ!���"�3�����M���˳_^�vuD��vy�4�vU��ʪ%�l)y#��V��N�+�����r��M��^H  LVv;���v��p�*ےj7{h�7�4��@7.bsH���������Wuh�+S7�M\Ox);s���w�ڐ6_����� �<�믰Uת�tc~�����*���rÚ����	;ʦ;�E��L�Q��W��oGPX�p����v���RY���Ⱥ���{{�H�C誌�y��Xf���eL�&2�6U�:���A+�:E8&z��[��Y�7r��G}�2#�Q�+r_�-��i��Ra�M�jk����Q�oq3�IN��jz(;bs��jN<t�E˰%������9��%������_�� nҊ�ݽ�@�3�ε}V'2Î�mT�37��̾�xtoC�ӥ]	��q���OLN��	7s�%��nK�:�9�>�����}�T��7������.Q�C$��k�3��i�.��{n��=�XFK�E��S{d��&�)�`N�ٸ��7�%d�˨yZ�W$�,�Lf3����[�Ewdu����:�f]8� 6a����ͤn02� �����腗>�2���cθPC�����;"R��5�qݗ�92���j�Z+jWs�2�7s�$�{+6s-�j�i7�\+���;D;��^o��+�9���}����v�t�Y�u[���ݮ�\��c��7Q��rs��Þhv^5`��Y7r�wT�����v�7��t�88TK�m�7��v�9��/ȡ���f)�̡y��˫�<�P��ֳ"�Xͽs�s��z����v�1��س�U̽�y�
3���W�r���eoM�i9��\�BH�PW������7M�ا���7j�˸���wܵ�9٪���h>4�\�b蹡ԼH�=G(�7��=�sC�)m�t�����F)L��Q���w���L��X5�v4d�^�|3u^���xg�9d[��u]"�r��Mc�1���د��߶��,O]��,��N��+�)��H�O2�v��	�v��ڱ\wܻx\�UUY3T]
��-�r�m䙎�ͻx�c�� 0+a�d��Q)��5���=G6)APHxaX�����=��G�R0�&�Ʃ��Ld�u({Km9�K��F��z/��;�fVmu�dP�= �ʫ�
ÝsO=
�l�V�ա�`�m��;!Uѡ;�cWa�!\� W�7î[�ꪦ@��*�{��}�X��UΉ�Ⱥ��fM=_^��~�GO�]7�����PjaY,�܍��[�M�#-=] ҮW��F��H�1�(N��/����\tjⲝ��!�k8���p��I�ɋ��a�vR�1V�~Ჴ����\�}v�v_	�Z�S`�n;�ҧ���zxe�B��u��j��0��LVXn���� ���D|W����9)U '��sj�����s�\��lґ�|syJ�\�H[uDO\�-���u�v���˩��ɣo��"/hW���N��N�������0:"&�����BÂ6�V��.�{&��q�]�E#d鎳�o�B�ɹuQj@��N؎"4^��W����}[����9���p�tӓ����MN��L=��ß:�XJ�r7���E�Q̙509)땚�MU�ٽ��=�½P��qgf̸�G���HXP�3�V�\TN��n��h�N�c��Q��S�`������qx��hV������gU����m��̇ >�U٬�ѝ|;w1"����v�n�	o�_��C�:>Ϡ�y�p��v����呥i�-5�u]M�M�ieXI�5�
�m����㦞 輌Ъ�U��	MԮ����MM8��M�B�_	-�(7xEM�-�p˝A�кn�b�c�*�\�ltL���P,£�
鸃rv�
nd�4��7'��Î�dU�ֱW`�MFN���\+,z�ڼ���9��2�t���Skl\ɥ�.M��2kle4��T���01:ة��s7�.�(s�/B���&,r{�vnr{co:�5�Z,Y���������݌˩ʺ�tj��f�"\��*��'E��z���0i�[��'��X�#�����jw���N�05S���3�ʋ�5�n�6/.,=��;f�Y�X굃�۝�	��5���X`wº�6�Bųӡ���s��5�(�H\ʙ�U��L��QNxw���ě��!5I��U�r�R�Y_n�߾U�6S��h��f��k�c�q�ʮ�ྺ�У��>X룧@=QQy4r�)��ӭ�ۑ�@/]WF7s�ZǹF�L�^�'CU�'ܥ�!�փ��u6:����]�ٵq�9�BҹwG*��(F�(���V��PF�����Bcv�pV�Q{�ֻ�kE�h��WG�p,n�����Y*糠5��>��Vf(����[ ����RAlwA��Nŝ݃���UnZ�����j�*Y[�`t�[��M]*�\j�D����
q���������;:'Q9ֻ�_�lfVK:֡VB�գL��̎�3&'�˞z����>�:c$�3���VVj�ǫz��Ȯ���!�g�!�X@ʙ�X��7��n\��h[��f����Wc��ޖk��\�5�ǋ���]vʽ����t�^W<O�2�b��f;����
˹��/M�ghI�Q��P���$Q�`�Ij	�q�!^n@���,Kp�-]Uswy§r󅷱W VVפ�9��̐;20�p=x0a���wf&Y��eU�mCw[8��e��o���\u�x\�DvX�9�tFJ���"�����#�闋�r3�t����[�Z�	(X�躋 ,/=�1�6�80���c���-m��a#��H��lXbnh[�,��r�U{L9�[�i^�����J��F�e��2�;�"�K67h!S*Ѱ��[|N�d������Nd)���U�/"NJ�8�ӌP��t�/W5���g� b�){�ܯ
]�����'�d��u�n6�<J�NuLa�̶'���خە�3x�]
Jb�6g�7��7��Ķ/j�.�ʅ��'BٛŹ:��^��T�Y������UãpKŎ�l[�0*��#y
��K���¦,�J�DF����J�H��ql^�zݸ/�;�g��i�ړ�&��l�h�����t�wuFC�a8�x���p!�*��R���-�tWt�	M���m9cY��u�ݍ�����W,rgc]Y�G"vq��Snx��܋�		�vf�D�R�N���Hx�EB��x_���79^t�B��0�q�Aqq��M+�N_]�M��:|���.����q���U��ns��v����joTZ����}x��f�{���h鶀9D�v&�/-�!��w��}�F�MDRS�}E�\uU�w*W{��OP�陸u*�ZS��q�|_RC!L݉���L1<�[���qyJ��}N�ֽЈ��§w��5w�8d93#�Uڑsq�F�b�>��ՠw"�j��Wv` �aO���3��|��,ܨ5<3��&pB����5Wc��þ��y���*�#;�5�
6sL�3=������įT����嚴,Wn�S���1�٪x�u���]�6�6(�_(�.+�g]����ةoz�#���8���\+A�o�v¹�ppB���Y�E��]���f�e����PޢG=�Kd� $�۹�g���k���ܭ����t\)�;��b�ơl���������jk�*�)-o����{����엢C�x��ϊWۋy�dˉ��KW�w6�v��i��q�yV���%[����� �
<or��q��b�ԗζD阤^
yp�n�H���Q1'T���u���#��`@vPad���K�WA^�|m�
p�(FĖ �փ�ᚨ�n�u�XKc.ē�{96ҠeԌý�.n�0���!,�7�$���n�Yp'�`��X�q1P��ub��u��I��<>�Ov���1�ԄѥVk�@��̰z��7��Y�;J��L��F#��c;9;�3��.Ъ\Н���u1�b��l�3=I����x�� v+Odӆ�3��Ω-LX��{�Ѳ���SJ7�ݡ�SS(�t��iڲ��o�/���K�#�l+Sݹ�G뙥b��G���@�o����Ț�ѝ�49"�A^3�Z�r��d��,�Ҭ,��x:�rv5X�������(��y�"���X��w��O	����$��{;G,��{e(.4��-k��:-VH�����˔/e���{�8�Շ,��s�ۑ4�W�1��ӻm�w1�(�y�)���G�v��4���L|r���N��jb�Gyo7���b�+����xWFQ���p�l�pv��{�YΚՙu&��{����"ޫ���/�:d�FM�uN���x%e;/�Ȧ�(7c\:��+TdX���v�h��v䕢����qb���43jƛ7�X��/�a�Fٮd���t{�o�֌â�-��ögQ�5�f�&��/vS䚚z�>�ӧ�@w]�;[�0 ެ����E(��񸊙AN�S۲5���
�sj���%L�U�سu�[����G����w�Sr!=�z��W�p���T��A����V�õ3�+<��V�[T���/��8-���Ta�L�ݴ-�]n#���S�`⎹�r��H:J�7�&���e҅�X�w��B���\WC�nc;s��[��������/{������.����8�J��LԞ��
dɵ�e��L;�Z4���U�J������ol�J��M`��_q����W�r��.�(��m�Y[�99�9Au��]�� �n��Oi���c�ݻ�n3&�:2*
���:�q���F'Ad�9ka�F,�L��ΧG�g�
���["��mt1a��ӑ������W%��sGP��3�s����s8y�#5�'!��Wp�뼛���J^��i��}��]�J�h�E��!����JR�jD�]\�@�=5��"z`�z���0ȧg��O�8���G�'��Z}5;�z���=/2g�RU���U�w��M���4�0VnT�1]�nS��Cn6�j�����|"�'0d���� �Et���	�����ږ&�v%+��<�Lv�E�E��ک:>��|D(�O��_|6oM߾#����-��BN�G���e�= ܁<U��Q���f�`�r�Ϋ�t�x#*�1.�ټ�ٛKT�Yp�]��������O�K�E���:�֛�k{���-���9V��a˝�`]�ON\�f�cPhuNГ�Om�Tk���)���æ4�9���
Y5N���s#�UUD�w��g>���Y�vrEk�C�b]�� ������b�1�fV����Lw�]3ˎKJ�>��{��L�3ڜ���A�wb�^(��+$,rf��N�һ�[�T��j��gdfT�B��U��R���b8�;w�J�^��\fN#���9�]�u�>�R����[���WN�9ܘ�$Wz�v�ל[J��'�2q_r��M_K9J��dvN�>2����s}*W�T�[����u����ѽ7�Y�^�Y���s�����]����t,�f�˵���y�(͆�:���%�U���ۅ�U�E��8��c��#ή�)�O��q˔��܌�-*�j�=k�ܑG�7)�o��K��X��_�Ay�}�3���K��4fo÷�#+울nZ�5��d�y��7��s�q��W=�����d�k63 <F4a���:��Kw&��Z�Ƚ����TrI�Ȟ�ȱ�����O}���'J��W�VRw�)ߵ���xv�������ǝbU�O�՗0c2�^�>}�5Y#�S���o�tu��
SF��@��;�6el�1k�SM�y۽���
�L�,�	ɞ����Q�w8s>\�(�˕;7�|��f�_O`tю�5�d]42�І�qq��uf�����\��|n'��-�w9�r�����}|7s�к��{�[�ְ�
^��5�g]��v�0��7Qz�4#�u�`�r�3�f.s^v!є�+`�,�U�sC�Y��$�E�7X��B��U�PŜS��8[1{��ܮ}��v�c�pLO,b�g̲S�/��	>������o:
W�4v���Y���嫋��r6nuKY��ݺL���������ǲ��~�3E�����m� ��kA(!|�F.���l�M1�vOo9�ё�l���L{{7�S�g�oY�����wQ�%^���5��R�U�`#VZ �����	+Wt�T����U��@Yu�� �;��1��Hw�-&�H�@:��B..-[��^W�1q�:ɞ�p��
�h=���zD��b\��rz����1cv�Lt^�ή�#*�S�f`o
�m����M���U���X�ur���qws�yBAJGr��έ�8��}�86V�6���6d���]�F`Ό�T v�*rz�'joo�怖��T��Q�/���!X�r��p@���Cݸ2F�F�*�*�L�ͽݻ\���׿u��m}�?v9�E:�Yu�t��Șnh="���3��;IuȆ�7N�ܽ��P���\H/0:`I�.�q����B;L��[�9Wp��S����K����v���ؽ��(���5����<2v�6���-���M|��ŋ!&��wR'�D��n(�-U�8�䜈躑�㢺%w*��ؘB�2E�4rc���l;UZ����:�R�v���&�e���'r��s6�օ�UZP\����F�ʸʸkdE�󛵦zM5P��6'.�/��{���f̍v�f.ا�:;`�g��<bx�.j��WA*j���f�b�cr�hnA����EI���z�P+:2礨�:㳱\)w feAţ���[B9]i�ł,<�=(\\]ӑ�SO�����V,�:��
3�!|�,��(�9+�W����(E��7����q�YzMw&vsw'�����vs��:�s��Ȟu�g:l+���ڹ�+���x(9���P��:��e�}PpÅF�M#R�q]|eP��Oq���k*\/�V3���p��ʼ+�*lOc�]q��G��1F{�)3u&Z�+�tT��Y�U�ވ�t��&k1�T�}���Mo��v؋/���ܟ�U��w�N����Fi�kf㘓=o��eŞ���5F�ގ��/;;;dKƢMOUw;Q2���$�\�b/��Ƕ�T)������Z��.j2��rލ�9jv���/���o%��-�Q�8t\�b��մv��rpÚ���&85��v%_v�
��RnVʼ&�	M�unB�0D����U����b��deZ	�˼8G)���Ӷ*V�;�+�՗2�l��C�始]6��]0��T^��ꦖQ{��n�����T��u%�q�t�X���4)i?,��b\����k�m6�/�n���ѫ� ��LoT�NM{#�b�-�ڰ��R�X���λ3�͘�K��
x`c/��<�R:!���c�xB�j�I+r2�^�`��f��Ns�`n�η�p1M�H��^ "i%�I�W��
�WQ5NM�Ƒ���B�,�}3�3;��Pښ�T\-�����ތ��s{8kB��]�����!�y�5�\��\6f
�Y<�a[3H�wٹ�C���m,��7UY�2���1|��xqN��]�[��[�neM`�g� �V��uF>B�)��v'��F��gTOo����=��H,�V�I���z>���U��#~����L�����赔�C���Cd8Q\a18����k�8��c'�f�S���s0��J�u��S��dL�7�t�����ѾN7I�O��d�>���4����|�}��[=��ݹ⣫�0�/�*T���O�*�&����6�?��O럮�H&b�^L|o�67ycw��2sJuW�{�����v3:��;�J�*j�]C�g�CQ'4R��v�;2y�#���>f�t^U����*�^Rɥ���6�j)N���T�]+t(����3�>�b
��*��ZlE���C�5SY����T�D�nd������4�6�tb��������BW�r���U%�'V+ҢR��I����-��8�{�БEL<��7<z���щw��O�C�{�:����Մ��	��un���W2va&��M�U���L���U͘���N�U�LTeV���O�T�k�<�����R�A�e&��[]�賂�PuGu�9ù��L;1�4�g�`�ˉ��b�rM��<�]�2���r�`U�ݪnr��-�-wb!�&�!1]�3D@���vEr�&F�'sy���f����b$Oۮ�+��G:��h�����}.G-�v���Qzn������7ژ5s������ϫ�`�k8JR&"��bł���2EE4�[J�ma�یp�I�0��TZ@��"b��[Kj�� �)����$
 �)�A�еIXQ�+R@+
"�B�44!T��8�JЂ�F-��H�����kE"����,D" �Ae[EX���UF6 �X(��8d)1bAJ��5�B�hHRQH�-!X)XVJ�T�
��k*�Q��*%T*,YZ�R��*��*�%HB&#��. (R��B��R,%IF
��� ��R(J�%m��1"Łe1KEU(b��B��R�eIY
 ��V�08n45�e[l��%&!M6�:� ;�;�x~�����r��}���`��� ��y��u������>���}�(w��=��g�9>�_X�0}�1��*ǻ�%��ü�����9�g$�7�{���gn����������ɱf�����㋂�ҳݧ�3�E�o�sN��l.���H�����7�t�k-��T>q�#,���B�-]�4�f�|���Ŗb��<�����"��	q8�  �h�8���n��Q��y<���3�²b.�)�=����HJ:����e��Ϻ[ ��h�1>TOQ]zd��a��H���1<N���\��p�@x�7��e%������0`�b"�/���=ڲ����;0�J�A���G����wxJ_�E�&@�0���<�LI@�7.�p�w�B�#*$�ɶm�rަ�d
i�8Ѡ˛Y�
�RO׷sMKY;o�J���m`�^��kBc���n�UDC0XB
lDsw���Ŋ�Z�_z�J]b?���cJ�;Q�5������+�9J��r����#�2[��n�p�,�Aw�ާ�W���Z��"c� �&ح���uU�5�0��\S�O1t{�y�(�_�k�nXV$��"���r7��ܻ[@��gP1�5����#��Ӻ�R0���/Ⱊ��ii¥r>JV'�}ȊSyP�	���sރ��ޚYN�v0cW�9��f�x�=Q�_7M��E��Į@��=	�W}����素�T�v�]�+"�m��y��U?�H@��_AiG~[���/XE .���R�z���\X�9��Y�m[ܸ8u��M��9��kQK����z9��������R*xdM�y��鎈�ރ2�6U�f�9aC�v9BӪ��H<ͽ�-��N^W,��땊:�)�>�����+�1�d"�a2Ϫ���'[�(���Yq��1���{��r}��_+ڀ���[���2� ��'.|�8��(3kM}�8�n�rJ
��?Nt4q�D���簕"�%r;��:��[��	��*|u?��e�=.-gɧ��"S����z�����w��8�8��h���cld9��q�J��a����R�)k����3[�G{��÷!Ь՝�7�n�h�<���mM�&�Y�XT�=��I��3d���K�|yŞ�Ғ�p���pM-6ښj� ����ur�\��T�"vyM��M�Cve:�ӴU�6�Î0'¾�[f�^�9=��7&�y(V�\zЕj���@s��cz�ÖO�p��
vJ�V!�2���� ⠲��M��斀��Ӽ ��`x���$|�0�I����k_1� ��t�����%	V3�u��9oRx���SV��4d���\�y���]��o	�L�[s65�O�{n�;(�%�u�srN�COS#����n��f�(�����2�8[����T�ˮ�G;8��Xj;�AW0[��ܙ���$�[�]��O'��>�t���҂�rц�e��Y�v����QMP����.�"R��֭�B���@�>���u��Y�%(2=7���Oڑ� �l{_��wl��m�b8� ���i��g��
^�:�>��t���8ٯݕ��MӾ�駍+���
���S���^t���|u��Ϥ��ό����F��y�m2�i�����3�\:���g�m��:��Վ	���[�Ǯţ~�{1o3��kޒ���d8�+���c��9ͻ��q�w�nkU��oǭw��������zO;�x�Įk_^[�[ɒ��]5��{v�յ2��$e�^C����Q�F,OM� �Ɖ��b�g�����|m>mϬ���|�(�^3OT�OWD��>�}z�=��������v<��H��k_О����X�Ҷ�@UL[ͪ�2��e6X14� v�<6��=�/��=gv��ϡ�>������_�v�_�}̻ם������8dT��R)�	�)FB���׼����qv��ӻ�<_y�����۟�O�H�	��L�d8���<��3����g�c[�=�B��i���H�'��������;P��&:[����_fO�TL*@<SZ���܄�j��~����}��9i��K���,��O�F�k���0EM���
H&�/ ����O�_�_�9?0�}������G߹ޤ �B�d���z����  ������Ҕ�/T�E�5͹�1 t�PK2Y3�|E���q���!����h��RoZFiy�K����w'�/�,fD.y��DU�w�q����״|O�<,37��+\:�Ȋ�8�c�HBT���<8A8t��'��L��%������g�4I��ְ�񽛿'n�k�"1)w�-�W��%�sy>\8g)�
.�Ҝ%4��W�2g��	�ە���� y>�B�Z!��Yx��kG+PF�02rRXp�Ib�h�W�:���&2���''�����&�Y���\iU�*7��8`�NĔi�
l7�n](U(%��xXB)$��39��8�XJ�~� �oa�,2�1�����MȜE ���5�� ���zb�����+�\/9����v2^�G����S�Um9!5�NJߙ�[�1������R���zi�<"f`��-=�8���Z�	TRu�
���K�}���y�>;����z
�k��y�Y{�,��*�������@���>�Ͼi��F��l�6��	�P�:Mç�c���қ���B{�k��6:*�8�DR��4/�ˁ=��N�j���p�U�f�g��P��pP�L����v��<�C�{8 f�<o175�L��C��yM�4	1��:gG�h���oxF�DÂ�X5*g6~�+5�si��K+O�x���T�x�Z4?;���w"E�MZ���s�Hh<���h5L=�j �>��� ƭ�V�1�Җ`�b�A�(�:=��è�C �)�G���Fȳ�9*Q��CB� M�I��[c���J�U�n���fƖ�zM��U��Ļ灌��R�ig��U�B�'��Y�F�l����r(��^��u��+��I��C�W��6�,��Y�v?�x���1l���U��[��x�Ψ�Z0a*\n㞉X*��V!0!�\��{�ܲ��0����B��u��iܒC!i�SH��W������`��݋	`�F�{ha����S���&���&<:�q/	g�8�Zu7k���u�'���~I���.yڇ��to��[������a�ԫ�}���`}��I��9����VW'0-!��{y�@zΔ�?B�֚�R��%���6c����b�Ġ�����7�"���ֶi�;�Cg2��rձ�*U
K�tr��mV�Ӗ��un��>�B���X����ͧ$���l	���0��b�(��Zr�WN�2�4[G_ـ�H���͠�}I�(�1M�{���[�L& ��]QUc�c6�lR�I<���J���w;E��^��y.�t�g�+�G�]g����=ϸ����:^=�Ym��\@�����	0Нo���g�׺<w�&W��������Jc�%�m5�=�����g3߆���N�]z�w/�X��������Wz�Lp��F�)t�mF5ڜm����6��t�7j����V�����v�uې���ͩ�ܽ��x�Z��x�1J��)z:m�ok�kΘ�Llw�:˶�m�yӗ�e�QY���-6���F�؅�8���&�o>nz:-f���$q�U����-l1�y�\�e����3jƈ�f�#n�@�<�M4N7��H�b���B.�[�\�c��r{b[ihG����M���*�~	�o��:���͍��Q岮4d�NQ�F�^W��o���f�OI�<V}]?���ϛ콯����ܼ7%�����C���Ӽ}.��A8V8������ `�a�-�USASX*z��Nzl8��}�F�� 7Sw`8��(���!�#^�d����	Vv�l�M�3�>��|����q�g��w��V�������j�=#���ti�7ʭ�L�g)�L�I5��񈭗j&�{J��|��d��F��-�vU��j��;gjiD�{-�ƕ���&�ƚ�u� �x�-k�zƏ����:X�Ufe�ۍpm7}qg��e�6�gҷ��%M�eL�4݆v�ͽ��NmM�7T��-.��E!�� �!�A��IQ�/�p�<���F̓��	�O��܇��~�����e�sp��v�3�}��u������x�9.3�|��;���}���9Q���j�VKE���j���VE�7��q��?6��<�lsfϤg��1A_�Y3/��qc�W��X޲KF�'6oۊ5��h[)xd�Ak�0�֍z� 7ì��f�jem�гґy_`���=m$ħQ��$Ť��h�K��7��I+$2x�]6_R�ΉE{;�Ţѓ"�a'�]l�����1	��X�\ҵ��Zƒ͌���cT������������*W��t`������Ý��\ٱ{����?.���WG��^�m�9ߙ�=���}gI�r�/��w�������K��r�����}��I�(�b�ǉ���aAaF@	�O���S����oګ���$d���]��'4�p�νX
�,���T�&DRc�3����ڑ!@����z��"����j�r����� �8�va��uS���W0e���>Z�X 0a�c��4�*?� 1��
T�]'������ޯ���-���?n��?�=��|W3߻��}PQy%BM��&Qn1��gK_�����5>�_x������ӯ޻�R�k����<�ǲl�s�m��roo��i��2�A�$�� �:���I�1�qs�.�5�Y�g�5�{��8���kq�$S�WR�_	G?��2��Aƭ:I/������<�+TH^�������?�qi�R��c��q��_�g�'b�[|E�fЪ��D�l��*�!�ۨ�#��%%��`��
V8���T$��eeX��Lr�}�ư�6"��(��i^9���Yi�4�e2�S9��D�E��ISk� �+��<"	X�X�"�a�+q��oh],��JUF#B#HSjɔ��]��2`��]Ȧ��ЊTmW�kQ�ME�+���M��JB2��
�
���t�-E�`�s����+��`!Nr�f@�o|8��s[0�$p�FMm����ki�6
K����5gm�l�܃��yoɈe�w���VP��d\�ƽ��mF}�f�ʠ������nq���ڦKdm�Y5#��ۭf�XЇ�K*]�/�T����V���d�E�Cͩ�(�+T,��w���.`�
L�W�$;ƶ$Ɖ�[*X�|G3lu��������x_��w#�(J�I���y�kZs�Zy���;�7�g�U�ɠP�vĜi�d#9Fm�Pf�7�z?�N��$eJQF�ǘ�D6�(K5��5U%"������3L
��uVe�Q{�N6��5�9�b��r乾�]���)EI�z�ѝ�b��?����hj;�\�?Lr��zUM��e{����B���f��j�iPF3�r��Wl��CJ�V�
�kN1�����V�8���p�NF��(**#��Z�N���c0�DFˤ��i�����ˇ�`?�x���0;��8���\��b�?v��ǘ|p����4'.;������f��W"���,f׌���ӝ�WP�1,ūbQ��Ml��׵�]",�z����JgU������-!�]�
�[W�TK<Jd
	R�$B"j�'+mV���zH�2#R�6;[mń� ���-����������P�!�!%G��
O}���{ɨ)S�˓��cA��]!Sr%�w>-�㵴�	���D���46�֘�J!�q�db�\ڸ�3iX$�9�ҙ�U��C�)��Nz��q�绪���$w���Y*��N��ءZ�|��`�Ѫ/��a�O���Л�w�<��>�����ΔZ���֎M."��qK���!TX#D��LX��S1�P�ޣ��D��	�����),sʜ΅�g*�p./��a��k�����7��mJ� ��bC+jX]$5hÍ���|J"�������^G׎t��tS��z����}���l�������g>a�;q��F4С]���h��-S@nԙ������E���ӛ���Z���L�, ���^8���L�?*��7@�.n]�ly����RH0��,1i��J	#0��jyQ[�I��c�d1@z<�"Ȩ�40Զ��$�{��AB;�*zhf(Vq�hy�W��R�
���]|Bbq�h�Fh�@�9���"J���+��-{��&Z$d����s:� ���a���Ґ����LD����-�VU��5HDTL���k��Y������0aaX! .)��E[ґ���Ը�=��YP��'���g��Ж�_B6Eɨ"g� 8H�*������-�8�*`���v�RBj������TVe@E`�Zi��|� K'Y	 e$ �3��7�oSP�pj4�ݹ�7ژ��yzs	��t�$7e�!��Qm�h��I�6�W>1n�h։bC�M��TPS�������B8͖�84t��9�ֳ�j�B��G"3��,�2��[�^��{w��vQbD3|��j�w�V�f�``I���)Ϝ
�BA'jR�IZ��fv����Z�djf���)�U�Td�÷�{��WZ�����
����3 ��t	�J��mf"�����-�p��1U�DB`�;Z�bDe���kq�/�<V ��`/q��N�VD���F�"" �,������w�۰��A���T!	E�5k׫��r,a[V�-��SZҙ�hH(m"
��b�O�m�B�0�L����l�gp2)QyTJf��"�>�A�>�1J��gz BK�J�;ij�)�7*�!�ɡ}��d��A�-84��Dsb���F��ƒԟl
xFʷ�h4L$����(�(Ҧ���B�"���dL��B�o���&�.�B@��ј�8�y� �`�HA�Y��I�ϩ��0h��9 ����`�}奪��v4w�-�o\�_��x{@�H@C`S���,�Y�`>B_~p"�����T�񹈄�54!	(ʤ�\�xR�[U5N6���DKc�=R[Ȟ�-��y�@��@� ܌�k@`�*���o=�h��"f�;���q$l����т�6��؜��ST��	�eZS,B\�/QM�o1�$�O��%�Qpmm<gސRT�mr�j�(�@�x0d����E�FH�PMYB�튈���lJ �1�(g綽���3Ud��о꽅�;*�00�i5dl���!R��ڈni:�j�%��$'���P�$	*��C &���:�KT�	DB�	�
���P��Y�{���
��BSűf!4�Nb�QWCg{l�� �)H��y�P�U��aFA��5�<�׹��PE��ǌӴ����D6DA�t ��.����J	�qG0V�Y3A@Brs��70���g��D	:�4f$�v|�3dJ��C�e�2У9
`gE �#�+K�PR4���T�P;�.n�"��vQN�Q��"1EY���0I��FGqX��9���BV/��`���K*�UMԹte�涋ʒP���#�AT�Д&�D�L�.ǼR�
����h�_W+{Q�҄���"hh���J��]<��B*��Nq�j�<�X�1T09l�"�*5��EdR�*#��a$�	�*VTwdG�Sv������8�+ȍ"(N2���22��eN �]��%6�_�¬�|TL�`�P!g��tf��wB�DC-)>��Z�*��	�!����]啦�L�Q"]�*Y���I)䇳�0�������̆6;�a�h�R�d�0h�ҋDf��1��t�DU�ŒD"��{_5�$t�5M�Xm%X"�RA�q�']!$͖`�.P��n�n�I;$�L^A��6�"�L�0J�!���|���1H(5+�%5)$�E��WT���2
jr�dV�ZR%j"P�e)B/Z��g��17�饐J���ݕox��q�~���r���V�Zh����o'�������E���"��vٛ�E7&$�7�n���j�zm	~7U��Q�l�L��X�h�/��"v������UM��{��Oj�-jq�������&U��X�Q%PBF4/�CqC	"
֏�%�"4�"f�vD��L�r� �f��b�f[<���T�ٔX�Rq��($b��\��s(�KҋT��j�,�����"$��)�3L��v�H{I�"�e7��]Q
&ƛ��/�ʡ�ز���U���1��a@�H<6�?X��d��;�ˉn֫��]L��UW���	C����"��Mf���,JL�\bb/�[��#��gL�@���):�`�U���Ô@L��[!n�-���^;R�I���c�&A�(}�v�q��E�VT
�	�u&���ti[X@�*ϕCө�8�"̎�4��xИ����NS�ɶ�L8*N
%�����MVvU��ت��C�>�'�6)p��"6�.��u�\6E�D��������8RR��͒(,h��T�jb�HB�M��D�D$��(�5t�)��>i�f�]Ew��G�2%2_��� D�E�њ7mꑝ�UT9�����O�_�j+����1m�J'Sm(�0��FZ*�&�*�¢�&�#��{�E�ok	���kR*bl���à*V�h��
�V@LR$��Y��Zި����-uK�h$	���UQsA�I��E��K�0B�f����F-��\$P�dLF LB3��q����...����̵4�FT�g�n(��
��g|6a3�R�}���1�R��O����҂`4�"��Yg@ج*w�iaCck��d��u$N4�+T�!�3�x�]r-\i�D�ܱ��^3%�os���V�� �Et��(�4�ѭ-�Jĥ�"�	������m<L�n]+]#��<uq����0T�y|;��*	HL�#yʔJ��Ϊގ�w\�no`������!S�o[��J��GV��b`�6�3�����J���b!�vãɲ����j!%�e,��+Z	GQR��
�>�;�����D��oŸ�$��RU ��)-#�DJ:���!��y��ƃ*h�P3�1��u�XO�E���XPXGG
��Qmv�>m��G�Q�*����_���57D(AM���祆��MPKZ� �'�,/�?�??��fZ��GY�0u~Z���-
�Uܗ1�LJ#|[&r����.�o)��<&�q���b�Z!��f�@��3����"�2z2������D[ڣ�d�$h�h�0��w L�F:�����{y৛A�L�Q9+
 ��H2����G�1���*# �b����������A�w���8�Q�����V�`��w��yjǜ)f�Ћ���A�������	*�QP�w}�ŧd�%hj�A�I-�ꔊ
�*��W
�ds&�:Z��B+X��l᭦4,�(�;�~M?�� 1�[:�p�_�O�| `Q��heLv�����3k��Dx$'�[���+;��`w�h�8GT[^��춠g�
�gSi�S�VA��IUI�;��25����p�0�̎�#8�)���C����,�H=�ǽ��╃�a�v-���`�)A4j�%
3*
��TgJ�ԛ}X9k��G��߼��
�S4�!�5릩��EI5U�mЭ%��h�C]LJ3�������*Jvx�6k3�X�L	�!j�jdE�<-�]���y��"���Dh!'�m�\�.-k��ą��94��T�egdAB�tw��t��^��3,�6�q���{I="P�j����f�
�p�#�"�q��b�Ү���䢪�HE븽�'���͒�4�A���$A��z���'
"��ƀ��;gL��$�YW_9aD`�X�lԌk5Dc)�x��n�0Y_h��j���Y��I1�Vq���t��E��e���	������ƻ�V�*艠� )���_	[g)���:A�H�";�i�-d��a#��8`*!v ���p�s��z���"�hĹ�he���D����1eA����XFD��`�
&�H��PP��� ���k�o`��r�
�|���AZ�dI3�0e}4FD�kG.��٣u��eQ.�T��O+D�.r/έ������L�9�d(.�H"��V��M��:H�T���er����{�+����h��a��(��N�v��w�'a�.���6��h�ԅ��^��qc�G�6�P_ �_-,60/�v[䍎m��J(��i�O151�H�N�GԄ\e�6�&��b�{10��+�8��������Fq�:�3qt�:h^{�*p�®�2�׵q5I"�J����M<�����QU�[���C���à���l�z�5��w���m�TV�#!j�=I� ��P#��`��b\�q�I�	Vg�ճ�xG\�/#a��(K�F.{_�L��;W�K���^K��p)rO��6��$5�&@�ǋ5)e6d4�הW��q��P׽�<����M���m2�c���|s�	��b(����YA���)lk3)�H���/i�څ���9�� '���7I�%Iڸ3/#�j��#mN0`���:�]���L	Il�6k��4�(V�Z;�$K{ƭ-2/|�
�ŰgC�7�)��ҹS�e�t��[�%Tșȴv���H��
���"B��Ңޯ�zM�l��rG�v��������q%Lp.�w۾���6��Xcd�� vA$���'T�� ����}o֣�m����PFI���dQ3,��;����m;R�|b_\WL��-��C����P"u &U+�3����<o�yР)�`rI��PS"��mj��+�qQ��XHu��@�bd9����vk�J�!/�2J�v=�vűTd�`��4A�5�ѳ��$�I)��,/#]I9h`R�B�Z��,�*6��1�<bC�B�K	Q����ڒ��0�D+�1i@���Lok�e,A7ݞ,�"�����;�mz�8^)�Q�6Q�-�,Y`F��/�������#�0AF7��:�n��Ȳ!�0�(�#�_J��8�D��Qj#	�$U���m�Q=���3�z�a�^4�عlaJ���U��X!�)�P�M�LAT%R��u�[���[z�k�(��=H+k]qm�'	 1W �D�jώL�蛌2k�0� ��b6����D	S���ȗ�@�"������֚h�\��K6�uں(�B B�U��'Og ����jU�Q޴$L�$ ���(�5*�h!"ɔ��$�A�PM���&�h�	4c(�t�M�:�ҚWNp�;�������#	�A,�!2�c���96��}3)�e�L2�c������#F�ю�:3�ӎE+�XިU+Z�"�;WD`<^�&oR�p2�)I�T2��DA��,�V�ķ�Bs�����&r`�!l`bQ ���@��LM��k>e�b�7��l�e�E�םL�KCBJg
rk��߼�Rq�
䠰]�W���:^Ϡ#\��`�d��La�׉s�9����L���̪�.�(�ڍS[b���0`P��	��[T��	����;ώd�O�7ȳ�}���K�BX�I$����`Bk�����,�H[�j�e>ҵDHS�0�sj�̢H��
���+۷���.R���Y�F͇BT�� (voJ���]K�W�|�Ƥ���Z�H4!�@�ۊ	�I��fa�1[+�yd-I_�� 7BFl�*B��v��]\nF���'g
0a��{[|�m�$�n�)'!����5�(L"I"����30���K��\��a(�t�^)�?��𕭥H�UR.�� Þ+�m!��C��$��8���77�����ȡs
`h�ޝ�	HRwd��lqͳ�Z�-FX���=�`,w�f�@I$����i�i'��&�F�V��)�H�E�E�	[+XK��%bP���z�j	�S�k--�z���X^�	7EQ�������s�$�d�7�H��$X�A
�-Pm[`Zu	�%И��_�"��cke���}��4h���i�����M�����Ш�D���X�����n���H�5.H! ����GCΕ���VȦ��C�)D	"hХ��~:��#6Q���`v-Mq;N��$
��<
�^}�b���2!6H3V
��2z:)%j+6H�PR$9�?!��
�d	DDC%�P�FFE��k�T�4rau)a� ���$�5]��$��8���T#@Ck�Y�q�	���h�br/#%u�� �C�	R����6���� D��T`M�����hLnRd�SP�pk1��fi)���٣K�
L�2A���� �`f��0L�[J��#�6R)u	`��) ��-�5�&���	U��+R�W�����F���b��E�z��q�>��T ��.�/IJ ��
��a��%��1@M��@�Q�{(-��>� ��P���~�����l��.&髶��$��ޤ(�h1%#"H�.H�w�\#�<p�L`��H$^���Iҵ:��H�!�fξ�bh�Z� !DT���2Aq(1&����9��]��2$k~)z�S%b	��f3��U��#ݴW�Dh�*@�2r�]چa ��f`2��E�ρz���B"
5݀�U�dk�ꔑ0,�(���� @�䔌W� zP�a2���ܙD1T"Q�������"��$�P��`���T �B�Qq&P��AaY�)eД�X0BQl�������
��(��5'��k���%��b �K ��h�6��p���f1��#�̀�!�"v��vzR�� $Y���/途� `f�����N��Y�@6#� �H�������w���Ę�gt��^v�9RWe�x��������j C�����Z� $���kaP�4H��F�U0�vE��pDE(�!��fA$tS����a"A��!��^9�ַ�� �HQ Sv	 ���ÉcC�n �T ��tX1jI�h���(PB�E��� �jԳu|U���Q�	T�B�H�L��vT��YBN�U�A4@�i$%�F��)�x�$��!
�8�^E.U�X�H(���QZ�f�b��eV
��Ff(ɧ��H:etq�ؘ�%�3X�h-(+�� �O�����$tt+X�"��H8��W%�c������&�h�
Ę�e����a48h!������cZX�	�]�,���*�Y֘���q��(�U	@V�h:Zm�i1Y�J^͡��2����DQ�����U��D��U�cQ�e�]X��W.�*��Uwe�c�Y��U]CA&Xa�9I�I�6�>�"#d��Wr���N�qHJ�6b/T��S4�o5�� Y�4�}gyL�ς���):��k�oD�*(jT��1#dI�EE�wjXD)З��QB�jYb�#���f�JAYh-���x�{h�`bQ	�°Nug�$�EB�(�����	B����PNh�����4H�D�g�P7+1)R�h"�1L�"���IYp�h�=Q$ݩ����=���������k�"+�������?�!p"��:�M1� ��8F�#Ea0�uz�~�t�UCJ�A��,l��.�ޣ�ͭGt�0�_7��i|׺� ��E6@�n2��2��f"F��n�!bd�B�<�k:����H#��\�Y1��+Wf��r�S���h��Y��.�9U}�ī��D�H�B�Z�2L嫐���0�c�َn5M�2(�da����%d&o%Y��&���'�>LJ���J�8#R;�R8���1��S W�ɠ!�`��uU�������N^4"�Udw6���mt�Lb��f+X��"^f��E�5CBhR��m5I�U�QW$I����k	R�QSY�*���-�X�kT���*E�{9ee6/�)O3�n��kho�/2�SM1�A���Y[6Q��$!��Rd�/0�H3��~G�6db?{��v�����?<��*!$"��og��V���J�MH���7Q�#�o����dK*mZTi�Xw�U���V���qĦ鲘a�)�7d�I�[U��I�� jQA�Q��H�;�JX�lTRэ�t�2e��ID�j�]�U��#W="�e"���EB�{�*n��I����K E*l��-er�56$)6LA�Z��E+�;x��Ջ��r-��dя��ߗ́��K>V�ŗ��y$�m:%%�Aİ��*��Y-`EA��ރ�g�IP��Ls�ZvPf�D�T�(󉜘)/m�{V��j��� ʖ� D{��}��`qsu5w�F�wR�7"��L�k:(k7
��zc�)�K��+޶���D��h6�����V"���!�-!�bH�v�����i��KX���]iگB\42�Ka�)��n��ќ��':��³5
K*!GF�wv��{Kk^�H\2`3q2�w���㭰\Q1�P)�%�ןW�|����@�а8琢���(�c�k������QDh�w`�azI�UH�=*,����	HQh&d�ZD�")���#���yW�.���BM��Ȗ�i4��X��Όm���ĠA5(PR���\!�����|����avSt%QJ9&�ڥfm�)b�I��F��g�������:������T�嘑�'"�vۜ[h��J�κ.b�������+{���	�1a�7�����V��K��]�E����@(6TR��:$�6���*�]��b��*�<h5��t�l]�b����턤��~|�Ad�y��)9�\�_��D&`0�����L����P�|'A3I�	@&h�B(��c�N��cb��cߛ"2���KP�HD��X��ZU0�X`4��)��� �����*I�L��+I��O�mJ�m@��@,d��Pi}�q^VgSrZ7�y!\���c���S�>?���b��AZ�dv��?#�ҕ����v�I�&Qwl.�}X������Ъ3�sZӻGcTME��A���<b#P®�A\T/���%hhQH&bn�R��w��³V[([;�q���d(���-�g�j�hԉΰ����ں�O%)!lX-�E+���k9��x�V[�uJr��Ө�V"��n'y
]�f��`��K&��}mE����0f
9p]B����@o6��`�*T����+�5��(V��r���L��vB-yɐ>uB��\Z��B-U��B*EU�FGAnu��3
��R�+܅q^k)�3��h�6�H��/������#8�,Z�Ăﺉ�KL)
`�*F���H�B�@^4�b&g�JFr��(��8B�RA�\�
��-KY��:��k�+I UP��{�<�B&���m4��
�2�E"PKƷ�b���Z)�%����˵S���*)�-�MbLSV�J#M	����XB��~���ҭj�"���h��-n"s*L�V]%I��Z������`�e|Z|?u��t]���=�%B�a��u��_���)�~=/#�9o!�����{���?�����/����޻��Ϣ1ߗހ�������C ?��)�%�?���{Q���Q��R�������_,�����&�Dw�"4�ڗ�-A�?�m�������3��Is[!Ƈ�|ߕ���Ti�n�˷��`�U��$P�G�(��	�~�:��u��&�������뮈C#�]�I�����߭�pdG�{���v���8ݶ�4r������=�D�$HMKJ�����mʧ"G�@v�����x��$�
PE57�ێ����}�MD���ʘ�D�������^��������O���`�?����i���������������3���s�@�%�Ki����7�6!�(' ��ӗ�Vp�H�������q �����L
�����~˸k�ic9�"O�O���?�?��u֛;�����!�P����W#����z"�k�+Jy��G:K}�.E\�쿓����c��I�O��p�K�qK��hbdh51U�~�?���C������gz����!CX[X�o:���
��g����z���O��� �!�bdS�Ȇ�0|���k�e4r&p4�����=gr�#�i�������EpB�8X�aF�(����H���P�,ګ�@0�����s�d��Fv����x]v�v�i�2�H��KJ�ʭ������s�|&��U����)�?�'ffE���p�ھ<ꎹOO�>��O�t�Q�`d|9��$�ދ�i=���[Zڦ���%��ٛ?躆����')r�҆O�sp&����6�6���?�2�!*���������4� �����i5����?>����z܎5�ވ"�A�⩠��{�[;�.`x�HR�[�r\g�ik���O���r������oNz����}�ʩ�]��N��͘����}��&�!eQ)A=� >ȿl�sJ�:�͕�]�C�;$^_���]��q�u�t�f�������蠝O����v�<����	��`8�=��9"��?���Y�{�m ��E2^�%6s=�(ρ~����όϠ�AT�'�|9T���Dz��N�q���đR,@!B(�^U�x�23��������(��;�q_'��^�ގ��:���?�0k�(�$��� 6'�b(��7����?'��#ꓹ?Ar��x;�oO@��@�J]V��~<�|Ns�o�;�r�rH=��U?;� �D3�G��ٖ�o�?��o�{�l5ʺ.�˳����1��^2�7|��i�ٱ��[�;�P~��?9TTSu�r��>�d��M���O�}��=lGfC5"؇�/�~Pe�<6��4�B@t �#�f^� cIT^G���y�:u������3����G�s�Ix���j�a��?��Nz*��fLDUi�	��؃a:~gΩ�5�6��P }ѐ05KM4�E�����
���U%Q
�TJ����A��ŌV�E��Rє��j6����KT�J��i
�E@�`�LIE"�TACUTUM R��R%D�P 1!MDR�!KHD�����S���Tyx�
1�Ym���JW�L�c�8��u*�ɴ�b�U��+Z[e��wiqQ�s���ź��uo�p Cg��I�eT���W��vQL��d�T� ��cv�`�Zm��J�|�z�&a�+���=����q���[Vۓu�_u�g\i}�����Zd���ݢ%����ou�R @�c��V�I��&*W8@}�0�W���+X*�IE6�b«5�Z�ci���aR��P0�2����$��@�E��y%�#Dm�jV��*��V
"�[e�*)mb��*E�EKj��61�)"t*#�e,��|�KJVU*�b���Z�UV�ҖʰV�DP�lAE*-�ĢV�*�V��F�
�")YQ�O�f�T[ZKi"��TTP*KiY*,��mi$LU��1�)iUQ�X�"�Q���ZU�Z�U��j6�+"�J
�*"����R�+mj�,P�UV�U�Z�((+[IUV���!����:��fWG����Z,c�f��u�:�hf�Kw�R�[Q˲k��mT�Du*�a��merW1l�M�����/�kTz�AR��g����/m4�e�����25�Y5mm�Tm(�¦�5J���fL�E����-^h����A��G5ݍ�մ\���]Jk�.�� C��)�J4m���M����b�`( �#<f�����!���
Z��7��*(��"

���S`@�e5V��t��G<n�6m�j���iJ�2
@)	%�#����PlE-�ʩZ[e*��aqb��Ŋ��;�>{�����S���N�XhuM����w}�[�|/ɇ5/�l�g0��lʟ����~���'������T�g��U	S�H=ݝ��n������!\�!���0�C�JAT����^�S]?e,߂�m��yͿ��~"{����$������_^�b	 �
   �$� dVcM]���u�[+2���Jqp1OXG�y8�x���c���?�?<z��* ������U�Kg�cpY:
�Ǜ���Я��Ԯ�A�>��4X�ƞ�@N�u�,���~�C����ⅴ����`}���$`ࡨ�@&ЀP���!$&`�Dz�C�D�v���[��13˩����
N�ͯ�V7C]���"��"ÿ��؇2>������6���uҚ�S�i5!�&�&}��@(&3I�T��� �HZi�DHQ����YR~�gpi�E7�O���dPT�!lN�@2�^E�Y�PC ���Fc��f1�C�a�?D���/��= �'u'�Т�%�gAɒa*E �I �#�(A��.�� ��(�����J?�?4��Ho��<~���|�C񎧛�+���X���dQ��'=?r�4+g~��z�&�P�H@��EH
�J�]�-=��=�Xx]]�}����h�F}�1'�bߕ�i�M>��B��IO��ܾ��/_�|�O���~��'A�'}�O%??��/?`���g�ɑ�1DT�0.�LF]�H��j#�Q��5;)�c{�ڗ���Ti��6���P�_?���ZC��C�b�Y�?Z��h�� ��ϟJ?�p:sK��P�i襭9Ԕ2��b�ȐP$!�
AC��@�L�!h %W)�� �h� xP��T�t���w�	}�O�K���̕����(��S���?���T��``X

�����~e�U�Wb�Te�:��:�L���8�*6��cNq�.�֔�Zj��n��Ɋg�.x�u�J���q$�õ����α��c�N���]���}L'�iB��e{�2h�}�M��)�'�h{����m�%��3>��%�����><���՝C�z��C�~ަ�ݝ5ױ�GS�_S�hXтA�545/Ry=œ�(}�.����Jy���#B��iA�'�	$��`�=��	$�?#Sb����J �n[��,���0l��͛�CMN2�C��0���T?�	?�G�km�V��o���,�vI;�"�T*�.[�0��g�l�>�֥��Dm�������$3&Jq��gB�+N\T�a+�+
�Y*b���P��E?
?ʨU��DF���jQJEA�����Ts���*���5IPMR8sО�W#6p�&���"*%�"d�s2���)W���%!K@I4��C��֌���FBa���K�YN9�Vj[08��V�W� w�(⠾����3�/����ZUSD�EV urB�9�'����ƖC�"V�PRQ@��q V%H����6�aEx���ˋ��]�|W1�f�IB:b�s�T�����1��q,EL�EQQ5E$E5CULH�D�E�44PTE4�Z5B���C� ��	�?��>��+��k�c�o;��̝�R��h��Z�Ļ��Z����GU:�����U'PԺeKey-�- A�����*�1�5?o�c�<��O�%ߣ��J�*�U���Z�7L }N3 �0����A�2̮�(�A��}A.���/���m%��aX@����vl�����əf/�p���������������o�����B��ߩM�W�#�;ld�:+���O8ە��'��$d~(���*5
.|$��(��:�U����������3:�X~��^<y[~K�z�����.Abά�$($�A%�5�Q�J�ʄTe����H@�be&a� T�b"P�C��`T ��E�fX�\��@Yo�$�V�>"��P#?�0����qY&���*%�[����k6��W0Є.D��R����R�-&�HՂP�˅2@Ml�Ub8�4Z�`���kZ�k��w^_ s=�B�r �!��<��ܧ��7��/�J%�ٛ�w�t�1�U2E��$>�/�i�<� �� ������o��t "l�{B�@�9!����v�V���� H���k��c�|n�hqG����UL!�a\�݀�>��G@��������B�mL�+��}E:h��R�;���x�_��m�m�g���x�!�K���h�!�85I�����9����"����og���m�)FC��*��*`PM�EG@������� ��//���U�I9����k�?s���М���{��~��P2'�d!�d��+o.%vC
��~7NBT[
�'�鞣���˟���M�aS�g��ݣL3u-��l�p���ZΊ�&vI.��s�O���D�	 &Dk����/ɜ��x%����s�C��o[��C�k��;�zOa�y���:��=w�1�&�����i�}o{��Ǡ������u�o�/����BO���V��8����R��&������D\Q���(R>'k�roq������:z�/ | ~� @@��� �/� ~@�pC�_���~Xy|����~�����H+�?�Y!WŦσ���E��/���?ps�Ӆ�MY��Y�����W��se�$z�9��D�&��G��U�����f7��r���2}O��}��J�N&P�3���g�h��z�X�n�//�C���k�M�^�?�L2�������.��� 7�?V��1ԯQ3W���de�Ə1�������}�ö쀦
B�&��N�a��H�i}B��1���%s�fiꋸ_8��Y�mS(~�}�tc�7_�C�lAI�=Z�ٳީ�y`�kNl����wxF*܅�ŻM~ޤT��f�d�OƩ��:�g�3��/�F����{�G��\?���I\^���[Xd�=O�\�r�N�[���]�^�Ǫ��\*���1ƍ��kI�]��AGs��>_\1/pG����/�{0yz����W{@��]ŀ=�w�?��{n�9>.?d:�pO�9 ��?�?��:`�"R"1��7%>ײp)��6��ǋO
�W��2u޵ ȋ��7����@�����ꋐ�u��\y���U�*1��N`0?�+�.�Q.�(e��c v�d��?}�mT��#�qY����ل��9�)�c��ʢH��$��-%QKMI�҉L�15EPٳfɵ�]��i(�P� $�y؟S��D[\bj$F*
#�F�W%c�GSkj�ۭ1*Q�K�ʭ�u���N�O�I" �$C�$� �z~Uˉ�k���ֆ8�O�����5N�Z�fQ�L9�mcM�e�N+$xϳ�䕤pw�wᄎ�}���a�vmj���(b�(�J
h� ��h�� W3��2�]21I9*�;$����SW��:K����C��$ �1]��5�����UC)Pы�0`��f��f��˿Ψ�[  `%��ƭ��7>7�)��5;n�;���K���uN���N(�9�iSF�CG�z-��O
�
� +�<%���Q9���W��p[;������x�'T�GW�Zڴu�����ޓ��~Hu���=G�����T�>����*/M�S�ڟ�=��T;����������r�����:Ǻ	{�W�(;_h�3�3�����h�t/�i^�i��h;|T�;��ͤ��b����x�7���LT�	E4�A��U��:K��*��G�D����<(R)�-B��v��+�L̑�������R�D)eb1b($F*�UQVЬQJ؊���"b����l�\�J��|i�^G�=��<�8��^��
�<>��{��PXrr�͜�����ş�ߨ����}���=U=�<�/C�(�P�(L	��h:Ӱ�����N�^�����]
�1�q�ƅ�dk&Hc6Dl�!� 	֡�К:�y��:�vZ����Ԏ2�����TN~��xMF[ho~\^�)�t�ϐ���rE�p{O^�|W�h�/�<J�/UY�컗�����x����le)�-8��!�]�B$�G�5E%C��G������T�'�8W�K�
���{��z��<��I<)�W�.SJ��wx}��	�Ov������f��~�N���������}��}9W���x|{��+���3��8gb�@�����U;�ME�{Gorw-O3��T��H�	࣊���;t�Ƽ#�� �7��ƗU��C>��Uz���)��!JP��P��4 �0�T�@f·�?���	�AAJAE*��8`L_P��*�ل����jgۃ�u�)Ԭ�^
SQǲ��{�:�p%Q]hΧ���N�����2����<���D�e�������>/y�*0�0b�7%��efaRˉw�B8�8#M�P�14�Qc3��Jm*�b�Q�m�������TYm��E��V�R(���QE�m(��5��T�l%bŊDA
f����b""�%Ѓ��n;���|��rW��x{�9���;�'j���R�S����e�L��v�q�CMBDPAQ]�y�x�Lo_�~�9����u}����_���,{�?��3��l~Og�ih�~?����ͳ���k�߈�/�c X��eG#�?��s�qD�@?��{�/�R�G	P%�t��,E/�}�@2zP�(3U�8�����5c�:�(Ʋɉ�n�Uu�����~µI�4I�y�8��
Ip��dm���JH�RDTͦ���?_�ԅ�;e�P�O�`B���~.Bq�*�X�e`��a�Y�?���|��/�*BP1o�r���}O�	q�#��}	އ���+������r��}b���y;)W|>����xS��}A/yO�.��O���=F8��əw�}5׆g�z������d�G/�� �+��鸐�QS:�;����p$<��x'y�7��Oc�-�7��G�\�G�����먛c�	�M�X��]cs���F~�ys\����v���%�t�I�gMQ5�8��﫡PgE�(r��EG�ML��A�x��o�'�|��ò���n<��뗛��{n��&?�^�p�Wc�%��r���t������������]�d�1b�a�dcXϥ�7ܓH3��Qe-
)�0z�Aw��P용]��[�q�\��;ì�0kQG*�긴�t.]�Q�d�ӵ$u��V�J��pHy��4m99]*�qd���up:��Nұv�<�����y�_�����S��O3��'Ϫhܑ	8�L ���vmwEH��O�W��A~�O��t�%{�T�E0I�?vp������d�I;�#����y)])ǹ�Qڶ��9\�vA�y��}s6�u|�O���l�����Λ 7�P�D�G���w�ͨs����݇8"R�j�����mj�Q;����x)X��Y\Qv���~���N�'�_�9������y�^�<Y��ǫ"�.��@��{�4ɦ`���;���?;��^=���H���_|��\��pIt��T�)*&���.����v˗��@��{mIWn:��������b��~�2�p��c�9h{Hf5CB���w5��t<0�A�Ȭ˜M�!�ʅ-4oY�����.}
���}�ޯ��^X��*hd���,��b;X�%���E<d:ʖ�מ\���!�O���r��w���)�z����� a 4� ��Q	4�5�������3�U���1ػ�?#�@f&�I;�Q[���,�h��x>�k�,ilq�c��;�{���t<���ݽ�\���œ����4w���sq_L��#��0�� ��)* �.�aK�W#������[ܾg���=�c;_�O5�'�K����>P��b�˄�L�K�Ӭ���Ķ(��hEG�8��쏸~�o�vv��ϙ�G�p#�C0�8!鎦��Oo�˹�մ�y׺w[�?�Σ�>��{�l`t��^�힭{�����p^�m���U9�������s|�į15����߇����G��/�N��|�0��qǁ���`^O����&�vz�2@�>�����ۿ:��T^�1|�>�!��)����U�0<<}���2��. uT������t��;��@sə5�Dp^�|n[u;�ܔ��6�[|��V{�}Q�)��W1���f��pr�����������t�b--Wo�>�ك������4ޗ7�I?0y���B�r�7,p�~o�Y�����c6FZjl$B�X���}<�`������sv�q_6����^�Ʀc@r� ��~{����%:U3kf��i�N�Ϣ�\�ɕF�G�cs֎�E_4M�8��4�������A�NĦ`�wԒ���G�O�a?��QQTDEG��A���}����P�ǽ��}�WD����C~�lO&�<�G�~C�y\�A�!O����������h��}��M3���;�@�ڛk,1w4�aU�c�1��a��)��~K~mJ�	�3��pxp�H��
zQ#�����3�:^�Y�?����"��p=H����7�\G�~h)��}'2��Z-���ѿ~��c�H�Nc�������2���q�v��H�A�W�o^zOv���ST�nz��_�ƃ��>w�����rGj����o�}$�7�P3Ƞ��
����%/�]�o��2�����",p�7��?�\`C^<gG���	U:��a3;��L�������b|瓨��P�_��=��,	�D��[�'1���Fuc���/�Fρ9%<.�U��IE�H��L�8r� ��}����{�:C��$���Ξo�"�2;�@9�O�?̹Ut�f�-��Ԯ_�}U�s�r�� ����>�A��.)�zP6����Y0A����
�f�Q,;����1�O��u!Pqd<.��v��N~'jj\��\	��mJ%�-��\�T����I�]�_���`q>���\s?���h�b-�/�a�/�3��J�� B�L���
����g6���'y�����7Q�췯E�����˲�o������y/O��n��n�����ӂ�_��:o9ڷ
�<	@�}~�����?w��������q{���ʏ���/����]��ݟ��?V��T�%$��F��vI������SpVe���+�vsTP`W4�����vD�P��?��3	�#�O��E��P
t'���T��s���p`�\/"�.I�!� s[���s��X~�QuĦ�m!�����E��rI����8�����Yo�)�u�5�=���g�쳈�����{����^sA�pw��& ����C��P�#��x��#���hX?�%��������GK�����K��_+���>�؛������N;�7���
!_�Qj
`�	C�@ð���������@G��(J�pϾ�}2��@h�Y���%�� B��!-��Fq�H��p���9 �f�5єXoH .̡���ҙD!�S�A�r ��w����Kt2U�SQ��T`�P�$� ܮUQ��o8��iWҖB!�)2E���Q�dV%�	mA��Q�-CEJ;O� �"��hg�P�ge�ɌҌ|�EM��g��ϳ쾧���;��{~�|7���7����O�u?W��]W��t{oc���s|��эK��' ��|����Q�l��O�1����"�%��/�X���A��(�6@�/���,�N��"���	�4<�BS�$�q��@@� � 6_c��y�Ok�o���]��f���u���g>m=P���P����~��>�'�����S�������x�٧Fe��i ����e���	�Em�aCU������15K�Kw�Eh�g���LղR��_�fD�ֈ�(�G���,c�@�`ZJc�� �"�%@�r$��&�/.@�dc���U�	�U$҉�N��]R���m��o� C�VCM06^A(c�{�+m�#3��D'҅��0��䋌(>��
=��
@��г'��w䔀[p�� ��S�>�?�����0����C�}?������7�_����������+�>��Y?���BS�Po� #��~g���a�S\/�-U $f�W�����i� ��G),���%[���N�Zi�!�<��X�X�Ӎd�!-���D"Im�m1�b׈����h׉b:&r\�#ؖ�.�QE�	��de@)C�[d*��B�h&��/���>�l@�7�qq��"����aTa<`U!&�s�0�����IV`��K�h��ń�@f@�Q0j,&���HGT�!�O���A � b��B ���� �|K��>b\~�����B��g��@���ƻC~A�bX�*�ɷ'�������<������3�A̹�$ȼ����Jo�<���`D'ȩ�
�ߗ�Ū�uG�9'��0�p>x�Z�p������h��!4'��(J�}E�X�����$5���Y��i�g#�A��闸�`�j�p��WT�-�ӋF�8��Ҁyu� ?�LAR`��[��_��<W]�ΗK���N���6���������.��j��܁���I�1���>zf������u�~"�	j�+L��>����d�z���QN;�~	��:Hb1l	�VrO�������9 ,�_��������>�d����*����Ȓ�	��x�z��k�O�����3���Y�Ļ߁#�̗�7�{��!�ǉ�#�cV���'�-�a ���K1F�Gw�����ɘ�+���d�����\a�J��iF�W W̭2���{�{���O����W���_��=����{��0�_���ړ�UERQ���&J��#ۮ�? ��i\�HA��%o�(RWw��Pw�5��q!��R�k!G����"C�w�=��x�XgTA)S�~�i��2�k���x�#)��A�
9�Th�?�=��{>��3�_}�-DC2�w�鈸{����T6�a�̯}���<�9U�!��$!�?K������!��Q�)�E�Ң�H��lUSf����M�A�:����j�ڕmdʚi��R�A�U�7��d�?���+,���ei[T6�l�� ЈlHW���ƯJgW(g�aQ² s�_{����%��E�q�ϩ�{�,���o�>o�y�9W�?����&�bb�L�I�j2��R�K�����"E(P%=�K�U�ꑪ�y���mJ������.�J�G�x+��,-CQ��MS+D�b2�����Ͼ�����3UF��:�����6I4��v{�3����SI�Fp�̦��h�5F�*�jL��E��Կx����j�Fհ���jʞ���m6��ڥ�)$��HB?�Ƣ�)j��5(�YKTKJ���Ԥ�����#���BI�俅�soq}ϛ����}�w�Gf�UE%
�P�����S.��	�se%D�p��-Đ�R����gg]Ώ�?�[]�N��lKkވ��_�ӗ1�`}���q�o��WM�V��ڠB�G9q��;P�VmdPGRq֦���V[)����Y��=
�^C����!Э��b6���wNhӊ���3"����xѩ�SWOSOWKKW$>pxs�"�TUă�hd5F�R�`԰������Z@ #�U��b�%n����Ƶ�\����"����x��I�����%L)H�F�EcL��BB�Ia�E���i��%S�Ћ�iEZ���H�J�֓D����֖bV����k�⨕\�?m`�'\�!xo~ޘ����}�G�_���t����Y����8����>zN��(��aEɽZ �C��B @� ��M   SE���РI�p�X�5\=NȦ�����|OKpy]�h����IuںVڦ5�����+��[��H�ȭ0)��k�S��-4����=���=��a���⒖��s�����f[oIk����me�9�+]�dy-�%��s�k�h������e��m����ީX��n5��һg6q��L2N�l_mV��&�df�-t��|�7��{c8��1�X�4[�6��l��p��o��-�Lsjɓy�m���~)�T!7!A&Si����G����bGh�ۓ�g�;�֠�#�Ge����tӃG��o)�}q��<α}ךg��1�Y�p�љ�Ү�z��>�������i�C۬h8ٕc�i��tژ�:pѠ�Ly�X��^�^�m��'7�i̵��=�D�;s&؎��׳�%���Җ��ih�e�vӇ�Qm5��'�-J[��7['m�e\��G�+aմ�Ulɼ��:�e�պ/^��v����\�������k�K\��L��\h\�br�5�{s���D�g�K��'�*���:i͕�ۚQZ:��<Ŏӷj%^��9;Kmz�^_�����y��S�(�ʫJJT�ɠ  ͧo+ֱ�M�_������5�=ײ�V����;2Sm���tw�y_���V�m}+׀���~Ӻy����=���ֺR���d��e�<<f��ڼ8מ�P�2ٟ3����t#�pMd�ǩ^�u�^]q�.s��>)ߣ�g��|i�jyӮY�N7���#��k�{O}|�j[��=���<�4�6k�aZ}�|6-�'J+^}�ݪ|��/1ۅ�.�-u�,�;z���.���;k�U15��Zk�^g���ь|Ӎ����۟ZI�iz߿=b�ۚz�u��k�Fx���mYF��Lh��w��º�)�jz�[<�+�2|y����z���I�~%�s����J)�5��Ϛ/6�N$׸�7�jG��^�kN6t�G�W�m<����^���6?��  � �B��ܨF�Y B`�����d�����"&)�*����
*���&ZJ���*ld�
J��"E2�-�����b  @�!Ͼڷ��=�\vN��r��\�H}V������ߦ��, s�@`�mƠ�+�$�b��F XL�Zʀ��1;�:7�Ҹ��̷.����h�j�;�]��⌣e���T�o�~��9�ߦ㶗�o���=韞z_Mk���Я15�ݻ���^�����v}���{2诎�<�oR��\�|�g�N=��v�b���}�k������*,�I}��}�m��g�}�M�Nu��^z{���N|G�8x��)�foa~�}�IW�������6�{��Ϟ�}E6lm?=��ďnmѷ��=�yǿ�ﮓ��1_���r#Ϥ]3�xB��
��[K�Ϙ�ꖓ���n.*b��nk�+,g�ϛ=g?��yM�N�p��oC�[�=�ٟ�7�5��礗�y���ٹK,}��/Ǜv��_>�ѷ��ooZ������8{|��)N6�����x�����޼{i����=�����[ֽ{{�Qj��2�v�L� ?��B����uA&�+kQѰ�k���8p��͖x�!�CPe"9E�ab@v��,#�*���%w�us!%ŉh�B4!Q�J".4f�r��<�E��豟�hh�
� �a����mBq�*\AB��>�
�儸�K X0�h� �VV!�$����4cm��省�@TB��c�2jaD)�����a�/�Xf�Ƕ�1h>��*/�s�
�m����a� �+	.4�p
 �6 �F�Bأ^0�QD�ɠ n(Y�{��~�W��S��}�W�.�{}=������}�x���œ���J#&�`�Í��:��<묚q�Ʋ���g���P�	G!e6��"�PyJ��a��ȖNU�I��!EQ�u�X���^�(�~�g}[����Y}�v��O�s�u:E�}�E�ļyN<	�͎�?k���n���{|z���v��k��{���+n�}S�<�����^Qx��.�uꋍ���|�K�Q63$Q����q�T�!a�������yr�ȟ y���ɂ�z7D���X�FS?샖E��KR@��������S��SO3"<����2��CE�YK���,�DB�<C`.�]����AbVG�t"%�Z�ɔ�Ek�!i�tiK�����	�+F���P�cxcDi����X>s�p�_t��b��6���:�0��r�v�j`��Z`ś �i�FE85�͕I'��G2��FI0`4�8P�7��A%�ig��=q�u�!��%��b�^P���beȉ��b����G�����-�"	�I�lQ|��I�ā�Xvg�H�|�X��.2�vHɂL�K<�ۈ�QR����D��BF4��,��ƕSKQbb�8�8��8(u�Й��
�҆�N�X`ɆD#4`�����&MiTDr"T���nR�	��%�I3p��4"�`6�2b!5Z,Q�s'\$�Q5�� H����t�̌fh��b9D����:l<��1���F�4i�������p��IA����ﶕ��~�]ϭ��m��Ec�@<@BC   = t�e� #m��?�j��E�pҮ�qB��t�R��3]�*�>�E�A/,���+4����k���R$�t�	&��(�&��Ć�hp�UM2���m��6D�f'�VW���lDR��2��%k
G)qv����P��Љӽ1�
��,���%���Vd�'!%��u%ťi=�Mh)�XHVS�AY#6z#.��>��)Z�8�a�Mrљ�$��Vx]�(Ji�*���Q�A(�*�: h"Y,�z �Б ��Nh�q1��"	�@��>J�L'̊�*�Μj�&t����R�rƨ�LN��B�L���L�e�(�,���{!<b������eS�f���c�]g�f!f�z!��AL�4�"�A�YQ�<���n"�.�i��������(�ʞk���9&�V�F2��KU����M��
�{�0���2�<`���u�=0�M$��㒼�(�����J,r� |Eh(!��@H@��+m�m�؉��+IR�6�ߔ�é�I1A��|�(h	��1��4��4��m��	��Td�j6j��&��9�Uya!*n�@�.��s�u
xCԺA+#�ow?m��g�+��Q�>����4Z��P��e1YF&�#A������~Wp�����
��yJ��鬱O ��-�����̾�#*�O�v�t�`^�m:(���|k�B�nc�lXʫ,˭���(���=�m�ޝ-��؞�ŉ�P �� :[%G�D(��P��X�s13J�5q��k���S�9��)Z����p{3�Iha�rn���#��
Iq��X��Ӑ,�O�0��)�ʈ�C���JCb%b�z�Kc�	1� B��bԝ:�U�?c��zOX����@�ْ�\tF�؇nˬThj1K���B�0��2U�*c\Cc�t�̠��Ej\��eTB=@KH�↍��(��1�n�K�O4�ʨ�\K��a/\)��,��y7��2�{�[0��-�Q����h�0���[��5�a6�g�܃<��Tr12m?pȠ�h��)�+�R8Oh"����&1)h��x�֪�a�L���Z�s"�ҲhF�K�`%Zt�M�ӴS1-4��H���<Ċ]B$_t�<�\�U�p�A*J��}C�b�8�ڑ���= �P���Zcޓ�&#�[r �M�HI�]v$��iJ�	%T�KC�,	�HaMl�W-Ta'�t�AP���y�t-50�!�Y8)�}ń�i�BÒ0Wr��� ��h�ĕXMؚ�	*hGa9#a�
&A�gR02$��>�6�j)V���k+�sj�6��-.��UB��� �y  @  @ '�����̣�Z `$Gk���������$��$l�{�F�E'� ����,~t��2!��T�ȵc�^O�,����n�^�â�	��u��j�,K�=�G�I�J��+h��1ɹ�@Q0����2�/�����@3�1NL�y��f�mq���'1�� =۳9�1�"�:I�B��������+�-0�Zi�4#`��d�8��q���1��>,'F��5%�>���4̹kf(��δ��b0e�BQ\�9�%D�5[9�V 
��<QL��3��D����I#�4����&���,B(��+<Y�������*�ęN�I]&$�^�Q;(��Z�ʻ�Q�,X�'�l�J��V�vL�|�qP+j��&5
ь�t��̓���p�ɍ a�܃%%���q"eDl���<V��3i�ZV7CCh�!���H(�b��
�PaܤJ^ͱ˜�<x��2#0*�.��΁�!��֪ۚ��W"�a�ξ5�A
QFz��7VprBu.�T�X�ʲ9[^��D�AxX��$��>2��85 �Bz�t�;����>�p�>0��ci��{�u�ʟ�� Kِ:��S0���c
��R�y�e���G�|�Ay(*eT�В���B'2�ضA�k��� ����X�ܐ��^�`_t�d�f�f�Xt�7[�����iS�S"
%�L�m��)��<F��*�9/S(ZݰJLֽl�|���CT��1i6K����'�3���rQ�	�-RGU�6Pb�)#L�����[���]����T�|�ˀ;�|�޸?w��.1��n�� y ^G� ���\��($�R7f�1������~Dg�8����s�V���NH�1��'�
�*�tY������95�&��7-�}�Õ�Q�HX� �9��H�T�js%B���&��`�ég5����o�R�#�#vS���;�a����rUaq+ǚ��m���9�Ժ������fv�3e��H���)\[e���)\ϑ�R�4X�l��&`���uS��f�Z��\[��AAe��~�1�ظ#��!�CZ��+�+%,^ &��Wb)U�UD�)NSOQE�1���"ꖬ��0���M�!��A:&TJ�@��u����嘫K8�<I��o��(���h�b���
��CJ��%�U���ޡ�x$LU篱#��I� �����@8o����녧�4㹉@�����E���a8�s�7��n1�,���Cq�=讁��r`��X
ˑ�$s�͞.�h�P�O�ZL[
dw��lHN߁/&(�^8��q���EN�0��Ӱ�Rax�HejfDeP6jHbj��M�Ჸb5�@tDe���5V��g��Ĵ8�󄎌�i�6T��\�G�%ȓ�;���qP�j5v�$����m'ZeE�(Q�\&k6se�%�v0ٓ�,�C�j��L�g೅�R���{GBa}i���$���IOl�:fM!�����m�΀IC�1����xq�q�9,tA�F,�C$cB��du�ht0�T�c ����+ �p���^�HE#T�v)��˜��d��ֹZ�9n�<Y���!��t�Q��"�����C>@  T@���z�ʠ�b���n�?�q���8��Xt����AE);Q.4�7M���Nr�h�[[J�R�����F��R+�GE�Y�	%IЂ��Ud"hZ�����ҙI�i�lN2���6A�@-��	!��&d���s�iV�ڍ��\i\�8�e�lQ�[$q�	s��*��[R�C5N2��Ģb(Di1�)EeT�	Ɣ��mJ�ZU�F��V�( �D��+�C�*l�̡�M��mT�Ci&��"�!��m�Q�"(\@&$T�q�	J�&X(�V��T@H�I��l!�mq�M��2�58�V�l-�N09�kj��ơ�
ض�IUa"��
�A`V�R� +	m	P���RAED iZP������"��	RTPQa 
ٙQH�D��]KaYu�-v���M�
g:�j��r
�ʂ��2�\U�CAd-
�*�"ZJ	�e1�4b�0�
E�2Bkd�$ESMP@ģEUPRD
P4�T!E	CTԕU"��U��PP�P���D--)@�!E1%E@5,	P��P���@PbD���b
�("i�� &���
B����(�eAUX�(�h���� ����hb��Ĵ-(RPAM%X��()ih%�u�/��|���=GQ�|��|����>b�f�쾧�?�+����6?K?k�?���>���/=����ڛ����������e~������S��+�u����y�;�㺟'�~��x�h���O����O��}���n_����gu���m���o���c���OR�B4�U5QT�ICLJ�%T�ԵP��T�E$RB�(�% ��B% �%+BR�!M)HR4P�Ҵ�SJ�#���
�@P*ҲAB�PP#UJ$B�+J4�QQT�@D%4�R""� Ҡ�H��RU��i�6��V�Ƃ���J)R�
ZX�&�d�2�l�ɵl���ڍ���R��Fě-���aV�F�[6�e��0A��lQSh"������F�h�Vīb��6
�M���mRFʍ��Fȣj+h��$&�i+aT6��e[#`M���Sh��Z
F�V%�������@���)(fPB��)
*�"�f�h"
"*�j�	�B �"�j�
����&�Q]��Ԧ�6�mE�F�[H���[-���ll��hm �I�6I�ڔ�$�A���dڨЩCJ�%*�H- R��� ��"Ѓ�Cb�F�mVЛB6��l؛R�V���ṾͪjlJl�cejM�l��6�+amm�3A�2/ן�$� U.yS# rE�����m���;�����>G�|�s�~h ��=���W�?[�W����m���W�#����'�e��3�����7������!�>������~����������G������/~�_�?7�|��ׯ���~G��ߋ�_����_�o�����S��~���\oƣ��#�>���M���������/�-�#��|o����?k������?�~G�]��_������5����������O���-����s���G��_+�}���v�-�>�k�=8
H��ӈz1D�f����	��Z��fi���j�����*"e��&��*���i������ �)�	��b
����()��������h�����h)�I�j��)�*��"fb��&(���"b��j�*jH"���b����	����"*�h&�����b(�h���*��
��(��i*j)���`���
JJ������( �* �*(�i�hhH��
�jhh�jh*(�b"�bJ�(j�b"��&��
b�����"�&�""�")����$����
"!�*d����(����($���J��ja�(f�*�"b�	��������B�("b���b��&�������h�
�����&*������*�)��(
�h&&����������)*(�"b"&��!�" ���Z�jb���*���j���b�	�j"���������������
*�����&��(�����(�������
(� �))�����b�i����&J)"����)&�j�H�*���h��&*����* � �)����*
*d��$��(�*�i�(��)(����������� � ����(��&��������j���&"�(�����"�&��(�*�a�*��jJ��
	b"�����"�������&"����
"(��(
�)����*F�&h&����"�A\d�(��_���w�?��ʟM�O�?���Q����T!_�'�~�������z������nއ����y��/��v����'v����������k��QP@C���S�0	����ã�?'�u����}����3�u����Ǭ��w����/��-�wu�}��o�O#��z��p?���/k�~��|F�/?ݾV��t_;�������>Sc�6\�l���?߶�/��8��ϱ�?������������h�^�_�3���?�����?��S�<�;�J'��o��� /f�#Be���+��;�D�C����9�V!����i�Q�����/39��S��~ �C*1'�'�7�xz!֐����&�%ab���"�=�Ƒ�5w\m�½�Yg}0���FȘ�jP����n	E�t��&��5��=�ؤMI�pYh%��"7|�$�It@|;�5����b����θ�8�4#�����x���
�<�T��#˨��t�9$M�O��0�a{��N�W�JJ*o7A:�'�����r��G�^uU��
7%WD&K���������\H�fv�y<�笐*G�^͉��̐֐nC���B��"nawc�6wAJ��Yn��El�PuعɈ��M�Ű�ق|�3�<��?V�R�[�+B�t[˓�%O#@�z�91�8���t��	�{Qsl��d�� j����x���P
6y,��	(˹ Í�TƪZ���uւ��m�~q%(�qP�g0��Mj�qD��5<24yW"�N�)��<��e��T������:��`��{�R����P�E�:ri�����K%�CJ(>a�������k��7	����m�A�F�bB��%�aIQ`~�1<�&$}x�`� $o3́[R��E��"���_�G=� ,No
e��A#�P�)�.�:Pf�"��fS�1�~n��e�^T��>z@�"��-a)s����E%bI�-�k^?%0�]�C��[�3�#�!��`	@�����%x5H�°ۜɢ9Q\ 3[v�A� D�%�48e���-Nۃ���h��R%^x��>x��b	V�����WR`߅�9pF�8��>�S����#�t��}�@S�g�RJ� ��~,
��V��S�He�>v:C3�?����B���I?�s/Ƿm�
�s�nR��N�aٗ:.r�@�KY�]I[O
P�RbW=���fJ�D����L��R~}d��P�?JB~?���C̒(
,�߃���O�9>D��~>��Fߧ�,W�|�T??���!��TP@<��B|��>HJ��Cȿ�|��*����I�<����L$R�!!�O 5(����9�hCV9WD'DZ0�����h́0_��C�U��!2q�P?FBV}�XJ�~��'�ɇ���� Q�O$Y<��O!�w�NL�'�a���j9y��u��P!+U�E)Ƥ��Uq���V�vd�l�O�u*G8�Vʠ�꫌�&ʥ)�I^5E�S���x��ҏ�q��ǋ������郮W�Qfd� m�P���� s
ɽ`s��껴�̝��a٤w��.�ZNYt�͌��Y(JD20P<�??�+ �2T����� �g�	���S��!�$.�H��g�d/�d�%ݪڝqΒ�ѱw2���P��pwgv�]�[9�����C�D���$'�Y�E�����+m��-�FAdX����)?�b��L��j+�V j����������������������������������üx�J�1��w�&�wr�֔( �J9V��  �
�`�>�`         �@  
   �    2      �                   c^��  `F     n�  @���U�F��             �M` p M�pi�� �,N    � 
 -�  8   *�v�@ ��4�((��AA@�     =  g]0Ol<     �  gP    
 : �&     �(PY��       ĥ)Syw�  �     �g�\     ���                                                    :   x     < �      c�ޤ��\ �     @�P   @� @ D� �(          @     
	 �R�  �(*���>
@��  E@
�(���R�g��7�q��R��U
Hh���� �(����`�      h |     ��`Q �;�  ��G44�
 �� }(�M�   D  �    (  ��TV      F�  �( ªx      �*B�@i�`�FƦ���G���d��O&�cS�j3LI�dL��ODm4�B4ɴĀ�=4�cʃSЀ  )�&Q�S�=4�O(�3z���i�h��<5O23S��6���4h��=G����Q��Q���Cj� j��$��M�z &L 12`�  M0C00 M0 1  �0& �  4<�)H"SLF��@2�     �   �   A�4�    �   ��)(�&F�ѦA�&����  ڀ   �    h           �B 4��&�L����FI�bbh4��4 4h�� jbz4i�i0OL&4h��L�@�A�?���̙?��,��O�ߦMߺ���v?oM&��]o�K��e���'��v�u�8y�|Η�x��$��[,Kg�;��l=*L�!��|��2�W���Y�-F�|�=���lNY�f-��K�o���>��g�5��:Wn�,7Z���{��I�\�)�S�\�K1���"N��2�D��BJHBϜ��,r�%��-{"c��$��Hxu8�BB@�z����It	�B2��g��n0����s�Fߗ8��klPj���t,�ğ����!'��B�D\J�, �#�HB0�O�-d�;i�u�ɠ@�M�6kF���˲�1-(��Y9��8�(� (��	�M`2H �$���!qB �`�PSXxaN��f3�uӴ�_*R���PG�����U�I����i�L4&�Z�ʈӭ�ƴ�n��`�a.�-<M�"8{ws���m��,U'1�D��cz���Jzۂ��e~��f�`K�)JUtD "����W,'$�[T�t��5Sɝ������UV�)�^��O��~�#�[���R���84�)��jMV��T�P	���\��qp�mbO�����w�F�|J�� �K�'�L@���>t�Ϗ]���Дp�)��/m�:��g���;�i���l�;.��l�5�~��Jh8h�K��T�I��L�J�EƊB@`�l _�!��%M��b�%f���@l-����vv7�M&�뭱�l�bz�7U��QRKTd��ׄz�Ȩ EP�=��Tp�`�z��I� �I���*��%�9��,�?)WD�����)5�����������x�`����c\dDu�F܄.(G�j�؊�!�/g�Q�צ�Uu�.��Q�Vg1!��?������r 1(\2'�{�P�{��S2�.��?O��p�*��-��=t�5��%��tM�J?Ga��i���f�R;}�*�D��]�i�~q�-'w[u�e�7���X( �
$ ��p��7w����
츩ІWBҽ���z��G_� �bA����DZ����0&[� 71��Si����"7V�ot ����X1�4ٔ=��7ח88n>�a�z,[4��O�k���zGb��3��������s�L�d�`�UH�Y�c�u)[���@������Jm��M������3��S]4F�k�ݒ�"@��&�B\A'��0��ݔ���W�<r����a)BRp0��ɣfU��Q��R��%���T���}��RF����[�#�&������\f#���:�p	G`Ka�M
��-�l����Т���k�������}Gg�)E�6��E)����*���h4�2��	PpD�?��}[�m�J1cٴH4�������2Hp Mb� �Lw�gg[4�_q�}/����_�	t	�*L+���?&i�R�^�\��F��޺&(""G�7g+�"U����W�	���ak:4��eq<X,7�~s�6�}->�X�2�X��	'�g�l@�,�L���a��9htM'�d��,ގq?z ߬d�	���>fa����G��\$�I��=D���b�����0)�ԃ�2��)h��j�ʺ��M_�Z(�IW=����6��m�H��+�R��~?j@��o�~�`z��R�q�t?�a��
u�ܜ�~� �L&� *�/�l*-��uz��j���~��uˑݯ�:�:"׶�����]����M�y�nժ���Y��BIHTUsq�XX�JR�ȅE0g*F �F,dC�܌F=N��4�j/tD.��/��8��[H�s�`� ��G�%�00��	b�$�5�������uu��u휿�ݙQm3�[�����vP�C��ٜ�&��\�R�G���M�JZ�����8�'̖��(EW¬��3�u����AF\��%��)�+�C��fQ3��0�hA���q��DJ#M� �}�֜of�G����}�!n���N�������Ͼ�j�9`y�nű�!�����{ts���>)${����y��A�b%It�7(�˓ę�_
9PaS��U��v�U9qr��v`�	#� �4�*(��Ɯ�[�A�`�xS�����!"�"o�ED�M3u�Ύ=�\�㟻kO�gd���\X��D�qS�}+���t'�Q�[ϙ�`��bL��d8�q�H0үug� �(tzdz3�FLn��uqF>�&=��h�h�)���1e�pb������|T����,����pSB�ڕ(��"n���C�K8�\(�,4�]��q�U�����9Fv���Tq�&��
����:��Z�������-���ʪ@����dsP{/%�*m7��N8�7��G���>��V�t�"�!�k-S����^ϝ)H�HfU4iM��k'u���KN��U��"p�8�՝�&���{�̳1q��U
Xm�C&g�.�FaPd�d�S�V�\�*�W�.�>^q�1h��L�S�rq5qnA����t�	0a����E���_:�/ǻs��[~�L,(&�!�b%2�	�f>RU�6m<��D�Pͩn-NoӜ����D��	����fWݻ+���¬3��A	�>�T��ma�Tn��=À�s������&�[\<dJB�%UU�PT^^���N��Q�� �{�*	�
�l�����a?<uDG�4]�	2f�}r�|�Ъ�d���Dّ�sɰi��_�� �6�	4"��(@EN�?
 �%7�f����c*�  k�G�p�d^�_Du˜�9�\��(*�0O>�� ���Vy��3ux�f��24��
�(R�QXi��'�jx8���Ñ��>�i�v]��{�]�R�G7q����gzs�����w-I�����?0b�@��E�L#�s���{C�{ �:���� 	�d:O'�o�Zdц�$���/�e�O�`��u'��4�~|66�i���O��Z)�|l�ݯ�
��q}<����wPpta11���l06ѱ�s�7�p6���>h�ю<|^���r���F������XU&�� <�|�y7���FIҬ!)�E�0���M�]������!�t)�h��I�O����D�7�F�8H	�����%.�_^���sD�
�'����d��aPYxA�L���r��i
�(ZGyG
!�:y���,c���e�m�N>�,���>"&��HlBb#{� U�
 ����NX��BP@0؁�D�G�Îa>9���'K�a-�, ��>}!َ����@�I>�!��@�tyК`��c��	Gs�e3�HQ��������V#���.�$���,2�93&:�	'�}�d.$��Z�Մ�ܔ�I bbbIg�"ed�K;��$�%J��80�Y� �.R���} `�'��C�����<y���N��޳^��W���^ ���� ��GF�[Bt(8uE�/ZE�!�'�| �)x ��l��8�>(�[J'��I
8�\*�.�J�T������Z.���7���ؠ��[���j��I�g�W����ݛ�GoF0�����<��A�w��o�5RiUW��Ez���X��ŋs?(��ߔg�_�V
)7�"=O2�*b	"0�K�ͷ�$l0���qDyR�λ�MTG��!JC|�" �J�LG�����,����s�1�V�{��5�����b|�{ Ҋ��f1*~{Es�}���"�m�Wa�1��QE���F,�#V{�h����������.���m��*�hR4ڍ��7�2���_��=�:��h�Ar�QH|�s1�X�46�4�]�K'�9*�^O�$�,�����+�=�=��
/G�I$�/�����=��n!X=Z��\мհ�*_,��f�`�}�EPf�E%b�)�$S��5�b.��0����I/>_	���6>��Z�>�50}�a�G�M|���]	���OTu�F'����dgeoMFSa�@g�̹< *��_�ӑ�_:�������m%���^���}�:�.>B�
�ga�����Y�	۟��ߙ����0�F#�Զ-��n�Ө�xi؃��k1��买Z�nS�N���A�.��o�@{�A�.�A)�b��5��_�&�\���sa{3������z����E|��g�Y����_-	�V�k>7V�*�����t1�e��T��ư���g���R_�Z��͌�{��'۫�c��mq[W�qQw9���s!T��_K;ϩ7G�^W|��{E�jYpX�bv�����f`������y �}��<�y�biQz,d�YP7�� N� �h�P�0)f��x���h%a�*+&52)$ƋEb�����=�ⴔHč�h��]hB��Jƨ�(ԑW�qn�6W��Y!$FIB$A�ɢ64c��U���j7}�}׉�w��+�޸�� �E	�H5�}���[A�����S`&N��M����%p���� A�,�(��ɏC!�:�hc�p�w��P�C* �B( AX��D" @�#`DX��R "�"�B*a1d�3��r*�Rr��N\���[�v���v�|�5����;l��F�Ģ BA$�32lk7a��s9L���! � )��q�*�3�if�~�**b�@B( ���(@�� A �H�B#�!�(�,+]dԇѪ�\@!�s�!�s�s��gBȳ�ozP��G~�Һ��Fn�s��\��
�j���o��� � ��ӻ����_��������{���?�����ቧ�'��E>����?��|ϻb�~���[��"�{��I���O������c�������a�_��_����䗳���ڟ�����_\�?��:�����Y�w���xᏢ�?g�v���=HP���~����ۊ�����'�?�b�)Cy���Q�}>��?��{/�+�}���������Nz���O�����_��|�s��W��/\J}���9KG����q�?��뽯�����[�oa�|�����3���J>�ߪ�q^��;����|��{�����\H|O�)h�<��H�_����^[����C�<���c��+�O���W��{qn��@U�����N�H�����]��������ﾔOE�����q�?`��z������oy�+�t��c�~��~�osW/����������>����_Q�����-3����O�z�.j�����p����V��_o��Ҵ����eE}�����?�T�޷OɁ���go���?�����/���~�����#�ȿ`�b���񽇷�>��z-��~��pzNkds����y[�z�ʝF�gUW�}�uw��V�`<���� )*���� ��ix�^B0H �A4}��G�i���8�����?�~uW����V�K��.p��'��m�nrΧ�f����E�Y�����8�8I�i���a��$���cN����mn���4!q�T�HTP~u�s����v�j�����!�nu�B�H�[�?��bZ�}?���]����Z ���v���-�8���9�� )���w+�ͱ�x���I_t�uH?�p�pw�����S�b��j��ޡ�@v~;�s�����m?e?o�Ʊ�ޖ�f-Z �2�:��C<�����;N�Y/ܭ�����|�����㷍{�8;�����w^<��	�G�˜� ����lӪo�0�kS��^��e��kT���?*y���x$��"��0�}�'��Q�~>���m7�g�9��uG�G9��0G;��^!����}|b-�(]ּ!��'�Fk���ts�#��� Lq��O���/���Bv]��FU
����s�s�ciz~l���g��gӝi��y�N;gp���{��*}h�����y�Ԍ��1���j�N֊����j�'����6ژ�_�P���3P��	�)_ɢ�f����M ��S�8w����>�6��}x �8<{P%�xlo�us�5��������+�?���v�p�}��σ����>ϔ�v�2�4zo�� s���pp�>��f�!���6�+�z�u^�/顝pٚ��ވ������ HppR���1�$��4��~2��?ew�.�����*}{�"]g�����O3�j�}S�G8}�=\�9��  ����?O��i�?n-��AO���[����s�����ke�<U���g�}����u������U� �~�����O~��� O�˷��������;C��9��L!����;Ju��� t`�;�w�эε��p�x{��P���I:�~��s��8u��_���Ż�9�&���oX/A������%{��o��C��cްa�éHHQ�sO.�p�z�����W��8��`�� G����N��)8��|N���z���#�
����� �l_ꓟ�R~�7�_�i��s� �V�V_w�����?4�@89"�Cy��s�uo�?wᾞ'��S�m�V_{�{���8~��M,b����2��.~��z}>/bI�5��k�mkE������Ç�9��:��w��~�O?~-z�G�N�}��8;X�5�j�q�|)�@�;׵s�ܩ���}N���=�$s�M%��x}{w���7��+���8^�zN��;O���������	���>��*�9�s�h���t>��Q_>+��A�&�z2D@}���w����8Dm�I�г�
+#�;���1z'\�][����g���rG�>�Ǘp�9��ps��>��#�~�Jz~���y׶�L<������#��a7�8 ��1ˤ>��i�8H_���Kaw6g���9��#�=��^����7�88Z]u~����� ���^f����tY�ڡ}SEv�z�}�K˩}*���z�ִ3�n{ 4 �888Z>%:T���ߎ���6$Y���H�K/�j��y���r�*O��~�L9�8VSGCmտ'nx�����Z�����oÕ�>﮿ ����K�A�Sx�"?G˝�ƿm_/%؏Ȃqk�@��  ������zS������)��O������]�s��A7��9��78;�o�$�9[�����v�������9«}V�������}���&s��N��(�B�3��W��r�M�s��	��7��|I��Ք���>�Y�����2�I�a_���',vps��
�(ctޙ�x�zs��;t���Y�c�?}��2���{�o���"�}+���s�_��{S����t����m\� �ŷ�ⴿr�$���}|s��O$KDO[Y[�/:��m!��??��8 ����|�88>�Rwl	�]5��5��Rc�6�={�*;��5j��>ڏ}��g�W�i�}��9�gCQVOka8{�n���������<L<��(<�⣇8 �|�#��!R�����%�☪�]��;�H�e���9���(ϊx+�F�����?�0U\��h��{���4���N����W�����B��'�Às���c��<~)K����9��?��̌m�Ï0=����vHpps����Oo��c~�"MG�/����Q? 8BJ��zl�5�9�p�_	M=i�H�ο�|V��o�Z=�=!�w�h|�6׍��k�����9��p���)��~����N{<H�H�� ��M~���4|t�l>ʹ��b������>�W÷r��_앍^�"�?�����/T��v7��'�yO��;��￶���6�?J�q,�܇ �6��8o?��:�{���p������;l��4��]�It���H��>�t6���8GZ�J��?N���o���Dx�:?�wpn��h�&c��������s�!����u�x�iG����tv�>Ǫ���x>��v���9�s������[��D�B���=��{
88 �3E�#F�??]�C~b�P#�N�����i@z�`�eI����u��q�I�a��8 ��� �c�?�~d�#?�w7xK���l|pg�?g���888 r�52*
)`Qf��˙*��K�VL*�'��ei���t��Sk�Ė*%��["��m%�u˻�e�w`MOJ�)�R�	��)%-s�Ζ�犸Ä˾��R3[[�S�\��J$�xJ��L��J @�P5���X	�)�i��)8���ө��]	HC �ܔ�[L���,�t����y��ξ8\�r��ɜ獺D����&���Z,|Su ʀ�陑l"��rX��E��f��x���\�Y��U��<��X�VZ�2ee��@օ�p�x�Z�鑡���6 �v���ݜN�JL���BJM�x�4�CU�M1�6��4,�+۳j�!�������<[8��(�-ok����^����!*���^��{�� .�z�4�&���CT�<�,�<��h�,�4�H����4�\�}v�eQ��jƜ2�Al��e���XbaG*0 �e	
DM8�ר�Vel���RQ�2�+I
�wv��Ը�$��76�u��BZj��Ù�ӝ#��-m�v]��E]!�4!�c}�a=�&�"հ�1'@�"嬚XJh�oIvٕQ+�;�5C*�f ��@����0 ]����F�+�Y�/]�#V��.nݗCa����D�YC\�wt�e6�h���ad�zI�n��<z�8���!:�qֆ���B�-�+��A#	��(]���Nր.P,׉HZ�رm��;e�(�c����Hr+a���b�I��G�%i'E�E����ݎ��0�DH����������e�n�٭��@�k�D�Cn�HoT�l!4�^�:��'��ٮ�`]�	s;v�%,Sr���P(*��e;hX�H�-BR�,��H� A�x��Q�-w]v���^m��}���k#�)7ir�9��r�ѝ�%L�I���	y�B�jgtyx�%8����!�)H�)jKL�!��Cm��ͺ�X���D��ܴ��	���h��M�"�q���VW#y�l�bK��Jg]���4�M��G�M'�l7`s���/;	;n��1"`��b :6Q��f�gYutN8��.Q#�Y4I��GI2����	�B,a�e�"i#�Լ��|Jǋ��bIb��1�!x�@�H��3sX�[�����\u�����M%45e��F.��U%��$���!�e'V ���Q�v� �c���`�Y�;{f����t���%`$`��D�WM�Q�����t�`�*-r�d!@�$��޺fѝm��Lɏ���u���o���bH�/W).�A��ڌ#yI�h1DLxJ��E����U��$��h�jW�4W!�N��4�+�E4ab*"N:��dw��!Y@��b\I8۴�Lj�01���ڜ�L��TMq'M�4���k���Z����^�g�Ygi[D4J����V`i(���pYM4�4�4���Ѭj3MM�k��m���E��p�D
@LQ�t��t��'qq
M��#����n����Nt�1	G]��ݚq1�$@'4��j=��i4��u�*��������Hb�2��q@$��ܕܯQ����*[�v�mR+	����fˎ	b�ݣ)�`���]���Ք�I�#D�i��{Z��׷bkJ��sMM��y�9��o!5�ݝ]�%(Nf�H�Y(�f΃8Ӎ����!�-��u�5��	/t;f�Yv:D�6�VA:�H&ܖ��hR
�#��8��qИ�a�������I��%"�#������.l�`� ���\f�NX]��B^P���R��R�vk/�ݻ����f�m�zCo\��5��nJ�I,Xuh�r����BBF��z�79��JG��G�wiM�`��k�$դ�.�0yf�0�ڇCV�!̳~d���<�RU$F�Hߓۿ6n�^�&Clg��&�����=&L�eH1e�2>)�'y����2I��;*�r�I�&I��6�e���T��HKB��]$,Z�Q6�"�*����*H�(^_��r�:�Њ�q6*֎D��ID�����=F��{��r�sҎl(�k$�Ȓ��ex����4��� D�	w�@���d�戻f$`=��qf���mU�[ @XkE��u�.i�RR��6�4���)�]���5��g-	m����u����.�Q�i�kBJ�� � Hh�#4���Z�)���˽e! �����S��gΔ7m��d68�I��j������|��g��8@��
ی�[Ja
A���+���^SGe��y��8JEt�q4���5&����RWY���8	�x�΋k8Ꜳ�Eŋ2(��I��9��Z��[���Ԅ�i��u��T�F��͵���%���i)�ig;�ibM%)��������Հ�{tvi�H�XE��8h�a��6�D&�y��:�bO��jb0��"K�L��gV$�Pا[�D�5�m��qM3P��6�mV����k����00����:�X��1�&��ҙQ	+�ɤ�, H����Gc�BǞ��d�	M5�S���
���J�
CG��$4�4","B�������3N2�Wm���V�n��!8wk\2����$OIUm���!ml�Ym2�Ik,_T�H`k��B֜:2r齥�m`�Y���2#�Z %a�nԄ�{^�5q�n���˝�	/;IK^iU#+n���v�k[2���;���ul C&�)'Kĥ:��6�"F @�Y�ݕ`�FN�٥"
�*�Q�up#���'���%���M�P�@Gu(Qiv�΍�k���Ou�M ���2 0)eb:��F��D3��[	`"�� `D"@X(B"B)#0�0`J�T�1
m� ��B(���P�D���D(��	�c�$�J�� J���RR}}۳�'�o�	MI{m	WV� �(���C�]bqQ�
�Sܐ�p9H2�Jfzu� �e����(��Y�͒��-��5I,)���v]v�a����ۤ	u��L��^)p��� @�{u"i;v[݉t�H��	���e����Wt#Y������g���5��V%�K�e3j�5�k���I��x&�����%�	m)�/2��-v�B��1,ݔAjީ8�� ������D�&�$�րQ�`B�\�f��D<���t��ݓՏ2;�y{���1p�Dʭ_1hM
2�S�wX�I��N��+#lJ0&ma�
b�,%���X���%�8�7�\&���晠㤵��d0!�[eA�cP��H���R]^����L����Nb�|͚d���l��/:q챠&Z�x�цOm��K�(�JdJ��0T$֙IL`�l��cSU��;6�������0 ��Y`bn����5k�F���ԻXEƶ��k��na��u��4�l$WKm�z�g<a���f��b4�N���#F�ZJ:�0'�e-�nֵ���Rm�4�זba�X%2$�����Ĥ�F��R28bz�졂&�k��7[�!b��Mf���p�I�%B��8�����v����m���v��1v�!H�*QݳL5���b]n�## BJ0���!��H���c�bכkl�h+�'#7����mo��q*2Z�M����,T撤�e��P����9e�up��3�WqN��a�jmsvʆ�"1;m��'1 #�Xŉ�Y\!��3K��%JW 4��d���9���k��[%�I ����Ig)�Vi�C��1�)��Xj�Wu�p����ͥu���j����`�a)`%�C� ���J�)�"ٮɤ jPi,�i*H�ke��E����HRv�IV���c|�q嬁:�=�i�5��tȚ�\�M J"J�*�(�k,�GU0�w[IlUc��) �d�nR\%)��`h��!	WV62�-�6�QW�!�]p��ې &�u��s% $+J@��yY�N��xr�H"`�2R�'6N�T�a+C�#�!�R�ě/19ډ2�T�l��b�t6�2� E� K/Wv�N�@��>���`�3�Y��,+%)V}^�_:�@$I8���&�ݷ�u�q+� 4�	@��[`R'lj�`h��5��z�HL%Y
���l��n�8d$@Leq,"���	_tݜ3���4�$<Ħz�j�e��\�w�VuIg6� đ�2���ŶR�X�!�XB�V��=�4�u��݁� �z�(��h�P0"ی��%,#�p@�(��IH.rj晠Ik��hz��G�e 0N��tċ`�t��[pI���6N�d8�0Wv[����Ȓ�"�.U ��I��XR@DH��͠�%Ǭݻ�d�!��������05L��`z��X�IŬ�J0y��xt�YN#�r��)<SW<KV,aE��BV M�ēX�UX���Κ푄T!��M�wK�Ǫ�W8` 6ˁ5�$�T����˱�^,��a:s��H���Z���	��K�t�n�q�9�L"�G4M6����
G}vSj��H�Y��C�-�@�T�LєP��!��G��$c*�"F�<�t u�3�u�+ c<ղ�]ڶ��v\�cbs'v�K��������K7t�! 
H	��@�ZRQ�s�4�Ě�"��e H3l9۶v����a�hA�[�:�GaB���.����KB��3L��i�62���J��c[�h� H���n�V2 ��R����M�+�aU2"���l����A�v��F<��H��� �M�D��iJ[d�������a�������'q������HbG5���l%Z+����5�nY��Ҹ�:�p�Z��AD)1�I��K�]�0� �)'$�E'	�gN�p��S�DC-�����b��[*&��7R V"3�@(����&@4���Q3M�md ��k�1#!�VH4Ⓤ�1��:���vRB�u�f���4��"B)���_ԁO��W\H�C��%S���R�3ht`H�pIE��ٵ�k�ue��P%�#�� �Lfi:�:�+@���@�B>%!�	:ָHb�v�4��Ĕ�)�Je������M�k,��8�B�í��GgV^��!M#�-Y�݇\�9L�g)� �9�[]��P[vn�Yݷ
�מ�.ipz��Mؼc"��\"α���p��� �kf�j`H����,dwl�0�)#��C]��$�A���v��H�wRT5�9��ݻ��zΆo�8�e��Ċ���̏�U�b�!V�\�%��8�^�]��q�� �	I�,U��{We��A��@��@�]8�H�n&,B�(%���	M�R�j+K�!,r(ɶ��I�|%d0�
[k
�,+'tf�:���<l�iF\��$p`�0�����ZN'n���M�V<0��#f���N終i�˨���2�"k�e��FB���3y�'����ᣪØ��Y5��XׯZj2��Q!�8�v�u���&٥���,��2�^���Գx�`M8�.l� �0'��v4����`�Bmlu��m��R�\�ih�H��J[�����`<�*v�6!r��F�X@��7Y�
�p� �m�9�u��D�Ͷ�nS4gM3`EQX@;Y��a)j�;u�5ۻ�ɤ��V������y�/���3��`�E�@e�.]PX�0H�8��4���[�����2r�Q3�n�W#��ۜr0�B,Nd�Į'wP�wc��4�^ݻ#�׋��	l��$d�"N�[e�,��bE�ԑr�Il`���%2��R&qL��CIjPdkjN�؉�@���3�a�&���z�@5�l��BQ9�k���y�v�������7��ep�ִ�U�Z�UX(��`���|5�(� ���
� �$�*BI,��- ���m��˝��띔��]F�UKD�2 ��{>?�z_����y?���׫�_��c����`O�3�D?���������QX����t�n���~��}O�u�q���kv����4�m�t6����H)F1ޢ��=�Si���~�}�'��^�eT�C��A����opa��,c�z��Ι"�H�U�k�Rm)k����	*���54�a8�4L}�M�].�~�m��V�v���M�V!"n�u�*����rI��Qq��~���8����&�}���-�1.���fL�*38�BsK��p�`�}7�@3��G�e�1�p5��%�ƻ�׭)+�?GJD~7��q���׽jELF�ܺ�`:�9Ů�Z�R���	�D�V�ښ�*�4���T���o:����� "�� %��I�+�i�8r�����q�%�ed�a%Y�s��4X��nG=O0�cz(8�����Um��!������'-X��h�m'N��Z;��y�4��Z#k��jj�! $��L����3�l�ș��*5�G!�4#ϔ�LZ��mOxx�48,�� ih��Rx�=��	���K@�3��R��J`���lXYJSX�ɮH��:}��`8;ˡ�
K\�5O��J
ˊI��*�x$��!�����ՠ'R����¤n��J��$��Tͽ1������� ����`]e˱<*ݱ�M#���M�%<f��K�p�2hy��F̂�I���d��HI��WE�6
GF-	~��9�9� �=��`��"�`��v�ds7�H��0F�Wݼ�BSh�K�
�V�
Ӹ�
Ń�>S$ӎ��I�]��9���6�+)�Сu'p��=��p���Nv�:�%�=l*�bn9��mđ"��X���/.:�@d!h.���j��%D� ��*�1�t�����'և3���p��N0œ���%p�:wf;n�S�B��@Tҷ�ugLmE�e�'%j�DM��&S�m�<9M*�Y�U���@��kE��-�<�Fc�3rt�Ƭ���L�Y(�1�T���*�Ғ�.�'��*�r� �
�H-���j��$O&�0OA琸XR�¥�$*D�����@ 6a�ѕvy��H�n�A�j�g��h"=gB��Y6`�P��`��t�����%������)`�P
��4Qm0�r���Qk�ԯ;R���:c�~1���~��Jz��m�GX��fN��iѤ��87���ӋK�]+Ht��-n�l`�U,��*5u�%pVU�������Ī4밌CM�Ԁ��u������Ź�M;7<����vM�<�E�k'r��Ά\Ó���\G�Њ� �1��\l�8�o�F��JWWӎ-Y1q+��Kd<��|߸^=���坻�^ݧ��j"�s�6�R�<j�<j�D,)6"�c�ko�>� hT�`Ŕ$i�Q�FIE	2 LT�H�Be��fI)��)��d��bI(H"Q�$�[��⥔Qdb�R���U[�%��P�U�CC�u���^�_�����2����n;�j����3;��oQ^w-M^ma�z_�ğ[���q�������L��C���R�;>�D�����J(��l3�&��
��������ՠ?����W�:����b��=��(i���{�_��&�A���`߻�$8��R=	�6�����L4�����5N�	�j�~�:���M�}��j����u�?s�V2�p/K���W5^��ؑk�:��H�@�:̕A�ۊ!ۚ�*���zSBW���/FR�97]���+m���Q��@I��|2)�l��O���,3�,��Jο��}�ݮ+#Ym�'��8m�8�'R�@�T��Q�z�c�U�B�m�	uhc�\0x/��i�KLR�s��q6�+��2j�f*e��ۭ� ]�z����A�5����P�u1�s�KM���
�*g!�Tnzϡ�iތ��0�5wM�d��Evw2*, �QX!/�^�`1(�c��H��(���f��|W*��bJ������m-a�dR��!��xzw��ZJ~S�#�Nq!ϓ�Q$ܢK�@��v� z;��5�/�n��*����.�S� ��;Ϳ�Gq�C��8���o�``Vp�,2D��Yx ����Dz���� ID=QuQ���������w�זC�����覌�A ��+`}�VʁdE���(M|�.�srG����|D���`)j	-��`�"k�$yw	�y�>�%Ua��维�K� ��x)r��s��M�?>�:�Z�|�˟.�۝2P�1ѹ��H_�U� ����ZcC�`�f�gsz��jĺ��'/��(�K�3�6z��3���f ʢf���\/"*�\g2�T|�A8�� �EPpW�=r�?h>n�ԁ� ܚ͕�&��(��-
Ӻ'/�C�: PM
�p��>�w4�@y�!�!C�<A���p#�6La�S�zQ5B��ig8QUJI�(N��c��U)gz��ǝ|,6!�{c<΃��J-���)�6"�.�L�B��pq�a��a�J�a�gzp�i,�8�׹�{���3X[�$c!s`M���{�ad��}ݺ�VvC$kexl<c� `]s4�ٖ`��4�4Ѱy�$�s�#D ���E�<Qj��}��?�J�uԀ�Lۦ{oQ�4=R*��x��3�L��n�j�aԞ����*M1��cT� s-��<A���BPV̽�PΜ�[�6`�	��-�Ⱦ��	J0��Q���ӫ�����r�����v��4��¶Y�9��]�I�~e��^�vG�K`���;m0��
����:x>����y��ß�3Ȅ0��/U#�f�0I*=�q'cXm�Md*{eƶ�B�!P%��31�&�����8�v�AEo�!�ڂ˿�
A�L��zx�����ZAQ��G��[[���5�����t�o`]�:aܨ��Q�S�R��
ǹ>[�p��=Pϑ��I|`�j�lA ��PkR>(EƂ���`(�e�r� 0P�"��2ߙD����,�����
="=����[����>�Jb���Ղ��="h�_ �{6�ؼ���k�K��5�`�\3|��J�oV��`ߟ��[�UO�_Ȭ�zr/[h�!�9��[�sW�ӷqHE�(,�$�Ta�;/� �����X8iUr��?'�\��Ʌ���v�̤I����ڃ1�I��م�^a�[l��ً��3�
m��`s�%K��/@�·�da2%��"���qci�K�
�촲�맠qF�[��ˡO8_�O����=?^�w��M=q����>  �$TUdT��1E@� ��}ۦ-��i�m&5js��f���!� �QDDd� �*) h����G�|LmQQ֩�ƒ���F��b��2�Z�Mta�I���)S��D�W�"'2 �B)�E���ɒ�XA�	B5��LF�%RA�!u_�{��k��7�{ڭ�j9�B�P*$��!�@�h�5�4e�r2�Ax@�*#ab*� �V*��t�F�-��8˱ʂ
	�i0H���d�29��UR1��"s�����(�;����z^k�9��݇��]���� ��	:%@qwZ(xmL�Q�f�j"��B��QEM+�IAh�B'@Sݠ%BA�ʾꫠH���,@��4��k��}���4�_�+�a��q*p�k "_��u��1���o�4��3���y����Iȇ}hϧ���s�jL���}O	��xl��T�	�'���wA߼v��es?���6�����
���@ A?N��h~�����3�ge��u�73��d��~�۝�M���-h#������I�p<_��������{���s���t�M�i�����4�f�c���Mt�y�b�\������ߌŸes|���>���7����k�ǫ�Ү�]w�ì��oY�_��r�"f��<P	�o�D�΁D���6�jq�@*
O�*�
����p0�@Td�E@B2@�"���"F2ZL�2D&6�G
��QVGb��R� ��H��7Q�j��WJ>a�YӢcB�9Q�iC8@<�g���$�Bh�� 
����L�5&����%�-�;6�X��Z���܌�)��5oP@��T���2Hi�T1�;I��c2�� �
��E<�"��C�(t_�!�]JՀ�Q�3@	�,�9� ��< �
:GIK�f���eV#d�d��
c>,�]�Tܪ����!��#h��XD@dP1I�RuqWmv�j�Q��Z5��#yvVE�_t�5�Y!�ƋZ6������݉�ԏ��Z�*��HU�TmUt���yVM_c�i�.���ҹ��@dYD-*u6�lҶ���i����mM4  _�D�A��P�GZK�� dVU%1�F����0"�&(�f2!kU��[%�76�ګ&�W5����dԟ�5�{M�[9����\���skj�L���Qj֋B# x�/:B���%��Y�%E���5����V��DdLq��F�! "���Z�lj�b��ERh���E�m��dڮ](�������-ؚ�XM�,ʊ�QU��k�̾7JJƢ�뵶��L��4		 +�K�V� 4��lK HaU"��(���UH �EUT�
PA�1A��$�Z�B���b	 �E@�T"$��@S��Add@D�@$I$FA �O�X"H�DVDRA	@l���y�����d�?�%���D�C��Mv�{�I>d�%i�d��[�Z�`H
&���k"L�r�r6�۞%>�%�Gt��dI��˼�����udI�&=�j�t|4�s��,�U�`d�3 8�"*�" � (,�(�*� �_�"�.�H��H�(�6�
  Z(�+mh�Z娭��\�m[���*ą,wY�|V�-�*$��Z�P �I*6�(Ԩ���+PU��5$QVDq@T-KF��5"4V�ܫQ���9�v���D�VL����32f{Y���bi'���Mq�=�p;��ؑs�ʑb�c�U�,-�I&��}�]�6�x���r�gv�kw�����:�WSZYaBh���;o^!Fx�% .�
�1�Xp��0��㦹�$$8�󛣤7Y�腏��a�q4�c�;��;H���,&땋��[y�s�٬�-���$��i� � Vrٯ�n���{��=�hQ�-��dX�BB����H֗>��'��)>��Fn�p �0e\�p ����I�E���2ӽw2x�_Y/y�-��2�dA:ڐ�����D���8:3��c�����6%�i��&�s^T�,D"����1f��˯��}z�L)�Qm�-���ٝ/�4�)�������%:���k4��aàOLw�XS<�`Huٲ�T}�Q_u����!���� ƪ��/[V�t�Ri&�����[,v{ssf��ȁѳ���u*�)�@��\Bҷ,;m�9t@̪�o�4dv�&f������c<���H�r�O<WX(��XJ���4����EL9��x�a)�����}�%��� �V2��`�l�� ��x��[�H{�x���!-���:�M�)R�.8��7��7��|ؘ�
�҈�ՅA��&+5f��4� B�{�Gǩ��wRk��-��c\ӎ3w��L���h�V�.�_2X{����� ���=f�c��S�wz�a͆���͚Nt�|ur�h0��\�����7.0��o=|�$wl��c^��9�U��R���e,��N�	Y������ M����,9�D"BmLIlr�c�`�������.�7tDw�pO��I�����Vq��(�2�RXk��O[m�A&�l��u2�k`��)  8�"��iz�Y�B���7��݆]��x�sωM� ���ғk�6N+g�*���k8LdX����6l%����L�9e��jM)te=U��M|�����bw�񧀞�Զ����A��n���%-_hܡ��j�ۮ��0��h���$0!ie�ݠ%�9�������=J���L�����R��#�x5�u�VBb�v�θ!�ֶ6w��3z��p0b�Ͳ�6Ь%"e7�Y�BV�8٫}e;4kDg6�YO���/X{J�����n�=t�HK��<Ia�f2Tց��׭��u�������{�w�U����u��8��7�ؒ�6�M���Y�݃�y	��8�|�)�bu������2�X0H����i�D�� e`� �Km�i:��ݔn��g� L�>���k��4`N�%�����zTl�gs�:<J�]�2��X��z��5�,g.k#���ē�A�_sS�b]4��ӭ��o�޶i�H�6�R=�6D��s�!R���l�[(c^f�uݒ�m0�A�OGL�oZJ�*�z�$d8<��g��'�4sT�$n�R{hv�ѳ�@�m��F�M�4��'W�tj�bBz-'["׉,���RI@��1%�7��;�,1<U՝��ͮ�ja<��nSb@0���zΨl1� *q�,�9w�'[���Y,"D]v��HQ�H�$DG��9C9�2�z�t��d��B�����N�יWh�@��0��8��`YM6��GCڑ� �66�L�u��lT�;���X��A�]޳d2Fpᓖ	$rȰŊ����x��V"VqCH�AtI�w��T������Fw���9-�]XtEe]Y�ۛ�y����wJ�l	�\��d}ցN�	  
3���ɤ��V#:�䱑�/���)(�Z��iwz�+'�W�$ �+�=Xl\X�dѱ`�a4V!/����JB	:��M�VN�SHp+\v�ݔ&�mˆ�I
��01W�%���N�=��j��B�S޲�w��H���d,�Z�n��_m�I���k�Ͻ<I˗GVq�wh@���t�]�d]�g�w�% 1ZG�0v�#���':\V���u'��x��hp���Y(R:�W!+�.��ܵw�Hygi��̥M���6�8CU�S�td��u���Ar�)��Mߧ��Nϗ��i~&�q4�8�̦e2dK��
��!q�7�*�dj%��j.kZ{�6ѭ^�k�y�sV-��u��y��\�5}-�-sZ+F�Uﮌ�D��F�-���8EB���������nj��m��+k鹪�k����Z��͹o��kR��F� ��]- C���|P�J�����Ww�}u�S��3Δ%�m�m��V�>��	������>��ɓ�+�hDHj�4*X�$�d�;kv��F�8aj�Q�R"D�R�M�ٜ�ܓN�2wp�w.�9wpQMvL߄��3ݛ�-k6���#&ɶI�bfa�8�!�RA(d�wv�cb܊�!$�!#!"U��$Tu���F���p��N�4wz�ʅ�}&�ׇn���7[����'g�:����[[�P�'���k���x�O���Z�����iwm/m��E�P}V��N?��O��ۗ��y_���}��6��Tv���K8��>7��Y��|S��!��Õ/\���>��:*��}�h��*f|�5���P�����`�pp�BѸ�?�������S��x=�����=��W�;Rk�?^�z��8[#���3l-�.��ӫ�."��]�F�d>G��w�{[>kOY�2��Z����jl�"z�y�#��ۣ��z⫊�ޕ��6�A�߿�,z���G���h�yn]��o���<�To����Ƿ��ڝ���ΤbC��;:�>�Z{�����X�]֧���������XE�mlD[۲󭩝aϏ����^=��V�|�j�҅�œ��ώ�����y����Jy率�h���;���>��)8W����GƝ�6>�/���1���7��<?;|/�;���z�5��W����G��U�<�%s?����[�n�_�[zz�^����j�������'~p{o��q�뷭���ae~��p�as�  ���.�J9�s@ܸ"��v��{9�8��o��	�.� *�`�"�� �� ���t�* EBI�Tm�mJ�Rط\�,!U
�  � A$I�T�@T��Q*H"(Ȣ�DU$ $T@@A-|��#$�"�8�
�j�耸�"ߗ�4z�\t'͛<$� q��.�������@	�*H�J�5X�nnd�b�Q�a
#!BLZ%7]΄ B�AR@�F�ێ(�]D)����U T H��R00Af�M�Jܶ�mS�]]�_g�I|sh�5����;��6�/���/��U�����"�.����k�s��Sy��k�K��W�{����Er2j�F�+� E�\��F��I&6.���B��7�륣DZM�� *� �[���R�\�Gwb�D�U���Fܹ¸}��yٹ�L�'8H3��E7:�ۈA�v��^�t�]�	��*�q8r�$�S�� ��AF(���X�Q4U���cy���	;�I�HLLb+��Wu�˹,КhEwWIC�� �)�{��� ��I(�Di5�ݾ6�R����.m-s��o1ww5�w���c��5��zX��!���t4w\�	�t��(
D{��`�'���فi�y҆F�j5Z�*���[��ر�4���<�)+sp�>;ow��k��(I&\���Hɜ�es�R.���|��2B�*>���xo��͖���=ǌ��?����}?��}g��x�G?z������{�����/�Y�?C�4�5#��W�!���W��6|�������%���Cmި6҈H��.�E	��W���[�����r1�5˟;�]9�0`���ru���9����%��fY����e���S-!s\��~.�(�F�
�*��؉-KP&�[]�T�#�����`D0��_Z����R?��n(0C%I"��%�y�ދfz*�=�8�돁�X����_��^E�E�e:�X/+�G���B�pB ?�2�Z���*\��At�gp��zd�� ��AoqR�)���$P)k��*_�<��]ؠ
K�����q>.�n���\���]�lww]�tXb��h	���0���q�ű^W6�9ش�*6�Z�洭us/8U9u����wk��$U!+�D�0$$ C]�^7����ܡ��2�JS�\�s�4�d��� � a� ��[��֍eŲ����9��ͳ�[�Ʃ:�@X������u�=D�����,�����=���@E�G|c�L���Q�?��{#:�OF��{�Y]�.���P���f�8�_3m���o�`m�Z�%NCNb�}%x�?u�\)ŔD�ӣ1�	-�߱�n�Pd%F�?���Q����r����h��_��Pc,�F�-N]4,�Bl�G��&	�X���A2�V�
3)]��"��A臨w,-�3*���y�DR�2�c6|��ۚMoQzy�Y��+ϋ�����>�e���8��w Ce:�MQ]�<��}н�򗨅b�o'I�9P�=���)��Nd���0~��蟜h��ߊ��.0����;���x��_�S�z���Q,����1�����
�9�ajp���s���#^��F�[*�v�DW.jTZ�z�ؔ�ǳ\6���Q�xH���$�<�Hn�ny���T'1Rq0�F��^d,�7;�Y��0Q Z�I^(C��������9�-���C~s˨]�vA�`7��L�W3x����_vF�����
+��]��}r-U"�GL#�������
c,gJ��G�#5�)C�8�cF5���]]���f)�$�+�S�G��G{+j�x�)��"'&��)�w_/�bBJ4^T����N�k~Zl���<K��s���( ����VI>o��5�:AZ�d��!{�72ˆ��x�O�s2���fʭ�@�����,Q�J��V�<��+	�o�`?_/kgE*�G��	sf�V�A��n]�NS�O�}�Xd����WO2ێ��Ty�F�}�r��	��T	L3WW��g|���y�4�v�ԓ�%�`�!��h:i��A%���J�Х�]k�$1Ln�A��~��9��F�4��WyO����(�H�)�Kx-H\3] x��]�^�<����AX(�r�5QsIӚ�3��%
R��AA�*IJx�2���Sv���r$3�S�.��ʦҕ3�<v�E)[�������t����B���$�D�u�/G�����M,��yЀJt�Qx���5�*�=p���v�nH�~H�-�xZ6�Z���To�luh'6{����2�Å�:;�O1��[M�\;|'��}�!%8�q+�>�N�q��D��
�Ju�P��*z
ٲ��PT��IO�Q'<�
�F�O���e���0R��lX�!��Jy�kUN8�CG�KZ��sy�t�yv�@�٫� D;���P��	s�s]yo�]�:4��KB��-��2Ѯ�Rh�NZ����a��#��=X��#�(;c�.>����.l��Z4�b�M�TQ���lc�;u�ak)�X�l��4���lGU�V{��د��=�.>�yǪ��&��i-�`ۧ�l����%0OΗ��L)�[NkW[���;x<�:ūxκ�=Dun�=��#!��m�-B�Ɣ0��XZ���)�=��R9ꅆ�`J����wz�ű�x�s�s�������f��0f�$#Q*R�TZ��!#�AP⠠@[/�t�d�c~z��1�:;�R1����O]����$�W��w1	B�'wF�۷��FܭȮnm�j��ƪ��KV�£I���;N�H �.��˺��7��9�cˑ+��8ww;K2��B�L�g�1��wXf/�b��s���^�r����R�knV�V�6�mWv������LȖ�fw��II ��0h2&I0h�Q�X�u����]�Ov�,_g]��QBFI$*QU�(���D�|뙾��-���d�:��p����;�D�LTB]�HR���Λ��m�(�э�`r��|[˗5�h�F��^��Wb�n��B�`0�H�$l�3��&�]���&��-=ו}ϝ���[�6�����^��y�/v��w���IC�ȑ���a		I	����x��<��� %�?L��Y���������D!�g����İ�2"!���N�i�[�Q���}���]_=^6�򵿴�h��}j��k��j'�j����:騆�0b$�|�Z~�۰��ms�8%	�詆� �]S �Z����"�ޚ����%Yk�$Ҙ,,m1[��x�.v��<���b�?��3���J`�B"Bd�I2��1��;��!#�rMG��k��*C�<��A\��,�� -�+=�{r�4p�`�ERI����ݧ��kH�.4��uc"��DP��_K#���ڂZ�qkR�*T�5�ρ�~��)��Ҙ^ $=!劕
��� ��'pC���
������*b`��[�6D����1K��jQ�k���'cG�3��h�P�QK7'G#,B�G�-�p�B�7~d�t��/�>�׍�q���^�n��{�M2�~���(�'NVZUR	�ai05,�H��hM��R.�AT� ��q{8���0��<d�*�JA�"b�U�8�9��a�\,i4A�蠵V՝C��Wb"T3I�	y�	���{9$�nDt�p��BT�3F�(`ñ��<�A�n;��:ΘR�`;�Q����Τ�)\q�HT*h�EX���!j�$JRP!�#ֳQHe?3�FK/�A�>�0I#?̂�t��Ҍ�H�_�2(�)r��4_@�3L
��_��'Dvфs�]���mX�]z$�)�#	�u�l.�hfa��-CQؔ*a&���Ewo�W�	6
�G���� �#6�U���8HkDc'D�g5�q*O�'�%��#$�;H9+��?'&�mG���N��E��m�n�	'EḱΠN�1�32�ش@R=��
���'xP��%b��wI����P���%^f�Y�Rqb^a��!�,�\�`�9��_;V� ��дH����f 4H�D�����`!�GmD�5���A91N�j�z�m��*�%9�5F��冟�*i��x���q5z8�#�!��$�G�~�L:P(ZV2p�W�|�b�Il�h�R	�)U�cC� s+ !$dEup���R��Ƞ2�Ȉ���!P u�7�n|j�"�wS{�Iyrc㬌f���&��^�D[�cs64ck��;U^k[��Ι�K����9�!���]f����wn�wuA��sm�X�i�Z-~b�y�\����y�NMbh_���RiHňش����v�Q[��ڈحE��}5W6���o��B���1��sI�wj
#��6ח�����sh�_MzX�_Nj�7�ε_	O.	�$_�3��cQ�&����Z����Z�־Ϸ�����&&��o���F����.(��-��1��;���}9�m�k�[|�Y"!1y�)=�61�S�sKlmo���[_krelb��n���U�;��������#V�梵�W+F�'��̔Q4[�﮷�Qk�_�)C�� 6MQ�TmƵi�]nZ"�ݮU���-�U�y�����k�slj戬��U�<�o-rص���P�aF؊�tBFIA./�l]$n���B��T�MT����f�(Т��3%�H`�JJ�#b�!��8�Q]tg�� �2H���H��mb�F��Z-����ꉭKj������u��+�Wƺ[��Mo�-�\�����B g�6�D��4��~�O�� �*;�˓�� �?:L3���o2x^�)�������?��y�_���OS��Xh�:y�+K�yB��:\�}_��5�i���-�s���5���nlɣu�1�"���1��Mh �j� !���g��+�����W;I��������o�
��aO��!��&OÎ#���?��	�����oP�P�:�7�/!����u-F�J�IO���¥K���V��;�mp��[��W]:���C��5���+sq�Z��8U�gu�F�t�\-�mr�6�kEF.Tt���5s���;���J\�r�*K�!3\廻s�;������V�r��ӝn;�j���f�BI���[����eb�c	���HA$Efg�H޶���5�F�Yj�sk�U�Z�˻	�����ͷ4U��.�-F���U͋E�﫶�1��(��mr�*��(�6���m�[\���k�1�_Kk�E�����o+�}^�@W�B�\��*��(鍿�s[[�W�j=-m��F�cÙ9�*��lb��m^mg�m}.�X�4Z)-�Q��*���X�m��׺�K��Ɗ�ngq��ۡi6�ű���lb�����Eky�($��,RF��
���V��wV}u�嶹����z�Ld!���)&l�1�,�M��E.��_ J�h�-CQ��aI>.��D�N�r"
�pJ@ԔF��j�m�_��
�̯��
|]�wuII��*57ح��Qj�mk�U��o��/tpE���h���Qd�]sb�1�VJ��kW*�"�&�|�vdܮ��[�mE����r�m͵ϊכ^X�|y�yV+�h�������slhH�Iwv9�&��6T�֤������H��	%^�����L�!wnA�1�;��ڍDU H��E� a��AD�"R%�a��*BFU%T)"�.�`�wq�ѯ��u�|[���"�7+E�����U\�n[WmgϜ����ӎ�bf@�� �K��I�[��K���t�Z�ӻ[����r�`�ڹ�[F��S�h��(�V��P��!s�����k��ww��wF����z�yxTU�"���m枻[��mnZ���m{^�ڹn�-�ͽݤ��Qd��o9;�D�wn˺�,W-�"Ƅ�/��[E$��ED]���E�,[��y���"�����B	���X�).�Ę��g+�(٥حsV��گ-�ԵwҾ5��h��˖�\�Ǜ�|k��5����zDw\iݵ�˅�w@ Y�F�К�mb@F�"EoT���Ԩ��-͝�1ngWY:�F�Dl��w44���$��r먌@���E%bI�P�"H�2|DJ,�.���z��dd�%@�K���0kr�iwnY�w#��B�>��5%DycʼՍ�k\���-�Q�e�iPZ"EQ��;�����d�͹j�;&\�Z}<�G97+�k��&�\�� ��RD��|PV�,S},j(���W�^X������+������^��s���-�=�w\�c��3]��Af�C'κU�>5�+�mU|� "��_�Y$[�t��E���ѷ.W.�{�yb4sǷE����uȆ�s�t!>;d1d����)�Bd�Dn�|�R@@�J������y^k^j���ڮ���Q������nd���
1�D�>w�����($Ѕݮ�L�/u҄�V<ֹѨ�"��-�$Ed�-]��9����&E�Ɨ�N��W�c�(�ĬI�k�p�E	�.���>ut^�9r)HF�*f]���(Li���!0���(�>�RB,�	Q�X���.ƻ�Hk��
+%�]��Hb�P��.pܺX��$��u�Bm��XLi��n��H��~�[��$L���n�����}+mъ6�E�F��J40�+��ۗH��j�cQ	U�\5!F����"�2B22 A_���;m�c��w����p�[�m߃����x����^�y/��?��?1�����p�n`��@�Ȥ�� |o��í�+��{9q0*����T���"d� �XB0Q" �|�w�6���l{?	��#�񚋾��_��7޳��Xߪ�g�������?��?Ɗ�����W-��>?��&�P*WuŢ���C��&oڥ%_Mt߉1�E��'Ѫ`��4�zV8��=韠C�	�f�B?���������g���k��?��������rxg-6bG�S��=7\�?�Ab{�1S�44� ��m��|�`_���H��J���灭�bX��*����li��D�w���hx8���� B�Jy�mn��P����0�
�5:Q(�9�~�J����g�t�'�7(/�#c9y�k3���(E���7Ԛ�h��V�q̍�n2nf�"�����|���W�����s�S��bj3��Uڟ�5�Ǫ�	�\��N�"�Y�ӌ��/R"x�����l�m�q`�=G\*��㽁t�{]��P�,��}^a��4@�4�d�꛼J����0�4�@�c�1x�<���I�8^���t�<��]"�Z��eK1�hh�����^�t�J�ѣ(�� �[|I�ú��E��WCwi�>��~>��Xf�p�d:���Q<��B�kCqr |D�R��iN��"���#�l�ʹÙ����|=9jl���γ�ΊX SP��KH呰�i�76.`�cj��
���K�����{L���[�y�g�q� _s,�iw�����U�5�5;V��v��{^#�(�*����|�Co��-�w��B�kY0g�˦�Z9N�wZ���R&L_3r~z�]-��ǉ��rQ-��a�}#��=�(�S�Y�c�-Rj����O;��>x��0WaV��NO��@a�j��i��*f�i��d"\n35�#uk��1�(%��=D�9C�hU��.Voӑ��7iM��wB�a3�:ZS^�E4Z�� &���_@=*M�pL򼖟�YC4̜&�9<�S�4�o��JT�8:+�w~�|���+,uk"�u�&�C�v�v]��C�W8�l�-��!�s��.b-J{FXĊw��j�Q^#?-k��A�k��2^,�b{�pp�:mV�F��᠉��j;�}"�<m��9�n�.�áL|���N���������:��Q3��B!�u�CS���o���� ��N�JϪ�'�;d�ϧ��]|22M�yjq�z��T��/��Ҕ�j:�����weɂ��{���"��=b���l���R�����+����QTuw��A���,�����L�QKh�T4p�DI���'e>�p�u}��n���GmcW`׍�_�M�Ƙ��]F5\����q�8j��4B���ѹsH�S_�B3��u+�9)�\�C��<����?`��:�ׄ�F�d�K� ���N�bܛ#��k��M/natf�FI	�VS+��d�x�C��(�c��:Ue+I5!�[��G�¿�M�1�ǓE6��Jf�sv����I�_x�x={vG�M�˵�Je)I�ue�\@�ڿ��<C�B.���hnߎ��[��Q�٤6$�LZ����U�=DN�I�7m�j7hI+���ȑ����<W�Zw.L�
��tQ�[��A�����3p�'La� (��z��"��p'~��uc^�p3�c��f��L��b�����x�γc�w��m�������2��x?��1}�.}⧊amr{�&��[7HJ�l��4��j)9����b�t�{S��IQ%���ѯǤ�D&.�������`O@  S���(��_�G�?���s�?��gs�s�8�����@_XW�O�T� ���_���'�!��O�0��>�U������%/�!�!O�e��Z	X���|?���%�M���V?�?Ƽ�?!�_��(o���;�Jc��Z}q��m����v�)���-:�eT���۸[#��9�9���є�`�r{���*�M���zX�,سq�[��v&����q��<d����b@�>�=�;9	�9��䘹��Vu8��7
DfKҷ_��Њc��Y$�C�b�x$Ti�b@k���NB����DjcU��I#àQa��T�YP��d�Q��N���H[_�0)΁�[8��H� ��*�Pz%^���DN ƻE ���D�*�B�CK��J_U��E=c�b�H��Qv\(nY^) 0��L�Ȏ��d��S�@F,E�L�����:S���n&�f��LTE��y'��ݐh���D�ʆS����l�ʚ�!VK
�H�p�e�Ӿ v`�e�&�1;�P*�@�c@(�bAä��AU)�q��(����do��^a���څ�N���R��`��hnc��Z�^nl�
�x��&�1( f$ۙ3NH����ͪ�^"Q�>�s�ܑ,� +�G��27��Iٽ\I8LH��#d�<���!��B�?D�i�-�j�o���c������#�� Oۖى��m�,���$�^ �0��P���h,��{�j�=�mӖ�h�6Sǈ��$�euhX-0*��9�W.��a�>�ÖDhF���m�o��"z� 8ܫ߁�������;Ϣ,a�^#Y�u�Ѫ ܖ�E��;��r�i"z���L �e'L�RH��o"m�f__PMp��Ù �仮N`]O�L�A�?��Q:�F�E�5[1+��j"�9jl����IG.�6�$e���"�Y�֕��4� ���̆���q�s
��I����O��GX��Z��
(�{�"o�9H4�bh��kČ8�
n���aJ�]Cj�y�}D��\�������� ���H"���*H�"H�$�zn�O���j���U�ݻ��}j�!",m� �$h��!$BD�$�$��U��\�EfZ��������%��f?^����o���F��2~�tZ�R�GP �|�;��ȏq/D�i�����-��A8��*��#$���lm��V+K.2hi%�QchԦ��F���_��n�"�ʵ~�Sj4m%DI�0����r�S(��*�Aj"X#���q���ok��;���r_s��yM���~W��x=���|������}���g��]�?���~c�
���OHa	��A~�ը��i4�]�E�$�&�a��eh �ƵZ�ڨ�H��"��(
H�"���
� ,����$�	"��
��J*�B"�R�J1	�T򾏪��S��5����<][�疯���_���=�/������ϸ�P��ʪ1$�s)�܇�����F��sG�= ��a��_Z�}�_x�ߏ2�}���[I8���� I|�A�ċ�P���^>?S��W�x��y��IK]��ٽ�6������cI�|%	NWb�PeV�L{H��EA�0=��!즃q��@L~���?�4�YQC�ٸL�uw�l!9)���oޝ�̓�5����>'Ⱥ`�ܹ�A�ݑ�a�]�Q[쫩�P��]|Q�vC���8��c����-m�O2�R�3�q���>u������n��bx��MB�3i��[�6\�D�L[���!i赇���)=�PP�~��LA��፰�(��x�R��S�k�	J ::w|�����5Z�Q�KԚn��!Q ��n<��G�y��˚���+�@ʰ72�ȅ��Lw�ؙ��e�������lDx�~�@��kŠ%���ir_@̊Z/Jg 䡦�J�]��.QO�T�CƊ|�+8p(K(R_�9���E��9?lgs<���4^��t�+u�s��BT�U��6��[�}�x6�Z�ؑ�mN,�8�2�J�;��y�4wF�QC�U��6��Z|���|M9�B>�E����/Y���R���ĺ�Ǘ���x]��(��]��� �����m���s��=\J�n�eO
�^ݪ�$�/�#��o#G&����tg�6�7;^}2Wb������g�q�`�Jϐ���a�*1�`�أ#>P���wwHOpkI2����!�x�?M^K=I��ymcu��8'u#m�B��粧��P,PD���_���u;Ku�)�k�DT�T�n����NG)�hn��Q�%E�c�p��3.�)��Rn��r��
P`!c\d'������K�ږ���S�J�����HuL�>��C�/%˻(iN�ʶ�N�|��r<��'��ؘӢ���&���@��|���P� ϼ.yc��}��=��@���\���-��B�*Pt�9bN,�줽$��00ܖeT�>��X�!|���t���*��0Jۃ���xa=�囥y,�0J�J��+f���,m<͜U
D���I�IhƠ,�%瞣��ՌAv\K�'84z�p��?J�h���B��^D���S�R6�����P�ŉ�z� ��5�!�b�ě{.�9�YoM���''�5��qa���R���hI�jՅ-���E�r�i��b
K�\h����r��(�����YՑ���~d��C�	8N��75�/rN�1��@��d]i�#�{!Q��M�Ҁ,Է�|�!&�j�l�ޚ�2v�Z�1cPr�45�4���aG�3v�V�'V/g,g�Dx�2��ʂ0�bW�S��ŭBsE��GB��T�nx��x\�Z͓P@g���۞Z{Q�`6�%������><\u�O~ԟ<b_"G���#[$O1@(U:P���B�=.��Q�1 �.QF\�Cp��mr+P��A��&_4 �u��1�p�d|Ɯ6��wJH�q�:�X�Ӻ�ݔ�ϗDw�+�Q��ۜm��"���6TwDK�qe5@/�p���b�y����M$0�Mϱ�[J�'5�\,F�}�r~�;&�vn$�Ũ��2ox'�/i���<v���[�EQ�}S��㶜#�EiAL��,�s�r�ZdДoi���B�V�jqh��[l,.V��]9���[�  ===O@z� O@ 
h�ۄ�T���
]�h?���3��|Yd�����}�Ј�^��A�}y��#������8I-B�+�����Y���%��?�{m:ޟӏ��vP�#�3mK��i����� �|j��G��3�dIO�LJ��Vi�څ��tZ��뮐�?��{O<Ï�z�uh����U�������Ǎ���Q8�fE�ݎ�� ���G��1� ��T���3R�F����Ʌ�䎮�l��	HxB���/�r�U+� ��JP�S~'dh(�dc#
�� DĔi ;��� P52�7T�bAk"��*x	��M4S�l��J#a�j��+=�28ׇQJWz������������W)�A�9��xH1��u�X2&�!#BFg�*I�A�Hу&U�o�H�
2�w�ZA1�L�AY���?Up�	>�u
ّ��C������c�H�g!�OP��Q]h[���%&���K��0�H�`!�13�!�D��Vh��!ՅQ褈	�a�:Ȓ� y�(M�! ��)�����MY��V��0,xB5Z��Y-8�q��e��+�P�4C>Z�/p���X�*jd[��B$ʹ�\c�vٓ']��3�q���ᐤ#����bYO��-7
gb�
���(f�4g�K��aA49����@;�������YiB����@��3ü�H�Rس��ndˏWz���y�މG��Vbc�<��+���2�P'8���B��˚�Q��	������ �%��V�cœ2(@DS.��GLJЈ�x�=T�Cz��]�/JNPZ�tV�1�0e�(�i �66a3[����c�!��,s�qߵ��z��b�
aT|x��mf��b�^9N ֜��Ck��M!JĢ%��tjL�9��v��0�q����!���i���ⶈ[wA1"Z� �t%Y1�WJ Y7�Dj���B+H�wm�I�6**��f@�Z5HDl�ߺlA-n����7��UW��wt�5�jTر�	-��ѴTlch�,X�C TZ�!`b"�!A�U�IH������������)��o��|���fØ�8���6�/�����G��?q�M@*��(���V
�
AQU)EF�b �Q��(	 "���)�)�x�S���|���e������_����?�*0?w ����`���WA�]rB8H����|mz�Q��U*�?o�==.�� ������Y<B|��G�������6�>S�d�h���y>�C�_�6��`'e��e��~�k������gʋf�	e#uR��oz��)��6<�=N�sr-�l��=V�i��8���r˂/�(E^v�<�Pyt(}-Wf�@~0�ٮ��'l��:t�j�5~����P��eN����[�3�@BѴ�j������J����W&��c��4ˉ��fJ}�۝����0F��[C�(�ּ��Pm��a�_\&��.��E�`G˲���K0����Rv*`䆢�Tި(pF�"@xo��)FRH�ޕӘ�i�����9A^�0��T��iש �/�pDJ�n���ǆ�������I3yGP2�Q�hKL�{�^[m‹k׸j-(�u_1�,�E²�Λ(Y<�T܎�+c���`)�(U|ƈ��#t*e�ٟ;�7���6d_)�]���$ʥ�����i� R𹆞/kQV^&���SL�،�o$�W'��%�&���rA�P�=�ơ�:#T�ai÷JѢ��I��l�����,Y�Z����+�-f�����d)�f�`�0��1F�c)�����0�c-=�O3@:w'�~�g�,�	���0(d�v�X����.3����j��߷*��}5�AԽ���C�uL�A.kt�$����St�Va�:��4*��8k=ή�.:j-ξQ�������Ü���X�4ڟ>���eCp��OJ�,-����_#�h�2k{�d��y����௟��t���$�A5���J���T���e�_Ҥ��CZr�;,4����qӥMU>-\ǐ8�f(^L�QH�z�l�`|�6,9�c�X(�U�5z�ٜ����ޔ���Z�[�����CL�Lh���U����1HR��.�ȣ��k�I��<�LCZ�gQ�V��(�D<���住��� ��L�f�{�L�^z~B�0��6DP�^���s%-ɦ܌�q\�;�/(x�Ut'+���n��+f���)��~]�.��^��]7��7�$K#U�8�a�K'$�ٚʐK�D"���E�5���7UM��B��/K�-|$�7.y�����Yt��x�"�-��\&��B��� ��7���ڻf��rۚe�R�s:|]�~6�����s�9]tN�KR�e��b�;Yɑ�u�0��6�=�_�|�L~�m'at+_7//�M��r�A����{�8!͗�u�qw���x"�*�i�4"�?T+
�:M�ֽ'��Z^�IQ5���SL����]�N��u]~��+*##+�.���=[�����Lo���/%r띻�X�ܫ6^� C;���s
�U�Q���h��y$�8]�)N�[��߆c�I�媄,�B�4�r�-M���F��v�=h�ۥ�� [a(ø���M����7F/��װ{E�MZ�*�����kv0f�uK����m  ��)�J�`�]�����ES�k\W_S8�����@fXݷ���D1�	�DՊ�F{̥(U�Vtؤ�&�hP��U�s�<�R��g�Q�$]6�4���yN��9����X�M��ݐ��*K瓘�|GG}i`���f >`T�r��`�s�Wq!�oع�ɘ��Ȏ��ˋ�=y+Z�[RK��I�[��U%�)�鰤�:r��dH��=���� � ��^�� H��1 $����x\�Ü�}����c�}�������4 *8���^�'�|o�XA�9&�W�pRD)���eD"w���P����{8�Xe�3�zns�YI��C�>@��Pr|�LQ7>�;2��Y"���������G8?�p�6��"�b��c+�a$T,0��P���db�r�lg}��~��<&g��P6h` �,q��Q V�~t��$�<"���� �u�B�=qLeK�c `�WZ���d�4SܕGV
"��p� ��ju�x(�e�R�P��H�K�KB8���C�Q��@�Fh��4w��Ѝ0[�t��6�c���M�!M�z��Y�0a���#�
�I�(�� �A��L DP
����Ol��P�:A@�H�0o�`fK^�ӵ ��֏n��j �P]�5�V �~1éQnhVLhql(П��I�_}���jX�3��%���+��Yi�l�W�=3M�i>�	
��R�&mY٭K9��X�5�x�PU�]M�C"��Pv���B%A.:L�!c W�6r�5�!�k$��`�C�p�c��;K�b@�A p�i�2����%�ڑi�1]e�̸)i�;�X�SI��)V�딥��e��� �JғL�R"�b9#-)\PPPf�O���E�8�@�Đ��Rb�!9C�5�j��5�Z��q��)0���$�ٙ)��X6�_�K�Y�zN��ƘUWB��Gyo؊
��	xA.4Q\�����:���#My���^C�t3�� �!tP!����2��h�ψq\u��R#Zq�/����zx��T&���=�.�ښ���ְ^}�`��AR�V�U�d�5X����5SL���6m�R�(آ5[ h6	
����5q�	 e�������F�W�y����n������Ok��������p�Sd
y#��$+�\!"�x���:��!�����5�x^o�pX�]��Η~��7Oxǯ�X���Kۤ7�}$�A�a�so�p� ;��`�K�To�\����ŉ�ؖ���D�
��� �����p������dA��f(~dk�'���Gh�,jJa�	k��W�|�,vM�>�c�rE o�H�.2���?D�֎"�6D�m��1\�s��+,X*DB�q���i�׆��LZ6k���Q<� @Fk1nt�+!P�$�V��lj/Г��ܼQݞ%�S��PEȗ��W�c+;8Ѫ
Xow���Q}��M{V�n��>k�43�pFy4)yBc�$�]\���|_�P�0�W��#��	KVG�d���y�?S��,�{~��hڮfF�˲�ʃfj�y�}�E��$�T���y�0�}0�z�쁅E3ΰ����'!�N�"���5�ZC#rЮ�;������1��d�)7��l{��_�Т�CN����.���"a�w��3͗:�|�Ӳ��v=�E.��RH�nN-�{5lq�����&p2D^85�����G�ˈt��y�Q�{�Dm�N��c���א�K�j���.RGWP�L���9l7�zq�ڊ7=����ɖ���UL=�߼5�Z\�f�f����("�M�PV�t	g��Q(D�H���H�h�g�˙J;��qof�,���/�Ap0dI�E�ޓ&U,�J����9�Л�eO�\k�)��I��*�X��8iҷ�c!?^��A5�񤁭��YE iap~״X��*R��I�w�d�A��L��2`��\�ڌ����5L�2��)�9?�+C�|��ʼu k��� <{Ikv�O>���=9`՞�)@�cZƊf[FNyr|?��<�x:��ck.Tn�&kQ�w�}S�ZA2�u�#`?�75>1�*�ɬ� u�j�hc�%�\�E��)�3��.�"vN@����L9blP��OD9�Fca=2�WqXun:[ӟX�9�C�.On��v[��6H� �}���4�#���o,�ĝ�Z����lG�����Zo<���CWh:dr�q偓�.�	i&fAf%	b|r��Q
B-�z���>y0JZ,�y�礓(�t�8��CX\!
P����YR�}*b]�2�JQ��:��-����8���8'��^1r��k�4W��4GX����9EO�6��B�2WM1�	��2x�q�K�j�Ȗ����I�٤��I�SOy�h~�¤-N��Hɧ3�u�	vSx/�s6cy���غ.'o'�=(�5�Ȟ(Qױ�j��L)EzX�BӍr:��r��84���=�E�+�B"(����Z��ҴҾx;�J0JnsW�uP�`�1�D3�-��%t%7�@��ֽ��"˃�i��֬Ǎ����<{`Eҽ@��U3��NX�.z�Jbس!�H��GrU�;�`g��"��P<d4��~֪��
1q�3WS���"��ܨW��+>t%+�u_*�E~,��e:?y���-+4�%҉��n�9`m� �X��+x�(p�W:� V�w:�>�E��]��Y��>��+�(�oA�2��ƌ����6�+�a2����!��[ܑ#���j��*�xH
?��6၍^
���
67E+�����'�۽:������4S|N��ŊP�[���F�%?'�A(ZZWN�}��<�0����t�s`�U�Xin+=uTaY�I�
�0� m"����- hZ���L���N���u�s��&i�]�ߨ�]�΅,ۓ�N�Q����=��@3�����������|ߔ��"a�����Q�>�C��f���D���Ô8�|_lq~��1�O��
�4��+�O�$2g�L�p�J�'�:d�9R��9V�%� ��_�A6z���>�g|���O����~�����W.�Y�?<ұI̒��:C�
h���'j��W� :�P�∩�+��Ϙ>|]�g��5�<zh.�������i������ZQ�o�騬z�??K^�;������YP~�#��bZ�gH�e�%$�
��]7E!q��"ed��)5�&�=�zB`9t�}� I�R0��3��̴̜�0�0`��M7��`aڐ E8���Ǽ���?<n6�{O��n(��m�Z��>�l8�{�B�0�i�SXP��t�d<F�rC��sQ�a����nuTy@�x�`6֘�	 ��AҋM�M	8��bÉ�
-D�����*��aE$�T�B����:SJ2P56SZDI!��)��ڨ�33��l��ih�j�,�>YH.����(�ء���{�N����H��*O�|Q�b�h��ޟ&�������2�6��&ꠒ�S
j s�8��U�L�1q)A�+����X�*�iL@O>��DM(a�@��Z:'녴�
�	q���$t	t��f�6���Y�%s�u��h�ǩ!P$Q(�)i��Q"�G�%�e�@c�m�BA�E(���y����NJ�]e`�Α���NI)�qrD,16)�FC�(uW�?��Ӽ>X%�v��;?�~��p\.����҉o"E(!$#��FH�XF�E� 8uBZ)#"$!&�*h`�ە�&�T�߲սں�l�u݊��wu`�PQ���Բ5�A���@�����x��u�ת���i��]���K��1�܃�_q����|�@  |�7���b)`��<}< ��,!J��1A�j\�n��zb���GcMm������wR��]�g�Q۞��S��C#��*�lʋٗQ��8L�FP]����#d�g�C���(m�'�}
���ڡ�\e��B�c8��ʵڣn08�ޟ��/��\m���6��㋴����NU-��H�U	ZZ7��D�=r�X�h7CM9�9��c��ll>��4ێe�M�8q�Q�E,���⬨���M]��,�׮X�wF:����9*ti�z�H1�WNGbsu<;x�q1�j���qO]���BFnr5s|�*��|'/
��T�U�י�9B�TOg],���2��,�aD�Yg#'j�GE^\����KG��Q�tB�޵\�m:����*g���sv!�p�.:"�9H��<�7������Q`@��]�7Dc$@��8���X4D�"�r-M6�ͫ9��������Ñ����v\�e��0�8��@cX�@v<�K��9,�O�����_[辻���nM��/Vq}R��?_��ீ�|�����m{��A��%�����1*	� ����! ��͎����\,��|��T|BW�����Y�=8��9&�n�!C�iQ��b���z��9qZ6���n�|~N���Xj6��1%��H��<A^���p�=늯^�2 UA�����K*J��P���~ʰ�I���
G��!iGԈ������� � 8δ=��R���J+�����yW`k�w�N�۸j�޷�rZ�)�:+�����ɻ��Ebj��_�}ryZ2m�빬j���ˀ��^w6�%��|��r����| �=H��YJuK����<�9>����<ԧc��K��dp�O�/���OP�����/�/��w��Cz	)Or�а�0޼�ܸ�\��.���������	�i� G�#Τ���e(\d���m�zf�}P�$vGByu6�9�N��L�Q�-R�����:Q��?����-��D˧}�:se.*��J���Io"����d�An���/8�o4��x�7Mp/[e��Gi\7�-R���U_U��'j�d�>6C�k�~��5Nڊ��S��Q�~<��.����_R��ί�F2]^8��̑>񍭸�r�y?m�^�a��!z���2�h�/�-����7�3����r�"փ�c�۩Q}<�����,�����ήy�����ӟК�{�	��nE���"�c�d�)Y���
�(��eۧ2��/�_4ﮞ���k/R2�)�9���{�Z4�h:�́&�\�腖���,��R�*	ּ�/{��{����)J�_E��Gr�XJP~C����Up�'�����z�|�2.�(D�2�NS3� ��KI�2�QgI��y�)��2�
m����0�n?.�N�x�{a��}p�WK�S}�jr8���f�oI�U�v��.�ʜ��ܰ��#��zKS�>krhJ�Ӎ<1W���(W�)�|�����1pO$��BO��ּ�M]�hźD��Ӻ�W4���6����#!�	��G�VQY��ΒN�z6�u$��⑿��y�g�=����i�6�[kgX#϶^��4� �S*AN?iN��[];1�C�-�u���q�;��������A���}�M$��6!���ffach;�>y�ƅ3�Cb�0�~)���H^N����3�v��� ��D��!����Cx� ܋��=$Sh�c�ɦ߮mKi�tT�N��H�M΃;�����<��e`�v*�N���Z��$��Ͻ�;c,��c���,�}e>��CDp#qq��>��f�f�~bWV���
�S���Ly㹬@��`(G��'�����H�b!�1L��0���ۖ�3ijHV8(-mI5_�Ý�]�xRmdPi���A�a+�ԛ��jy�䠹k�
������x��s�3Q�A�[,�d�º�$�E�����fЉ��KDэ�e�P���ۗ*�c�� wB�'_���>ѻ%��Ryq���$�1�@H.ўWy����A�}��D�:��-!�:����@�k�r��V���ð�N�Ύ�R0��-�eJ6oǐ.n�O.�K�7��D{
nVW1z=����u���d\�tIys���	ә�c�6	���u����^�:�8�Ǭ[�<�X:,�b��'W�85�t�=�/�u��wBW�*P@�� �L�æg���Ko��V�ۇI,,��4E�T5v� F[�'AibTN��!z��e(����ɲ=�2�)�&�	^���  k���=�~��[��𽠟A>�����ک����%�I ��R=e?m��k�x��﷏�����~���c�P߸�ۦ�z��{�7�����{O��K����������i�ߴ���/V���R������i��������j���}#t	�>:�����5��%�8��sD\R�Ic�e�vy�)�V)(�,��q6�(W��@�̠�!#B�Ҍ8'@~���R����a��4f�L�5&�����g���|C�s+���a�ѫ�������z����E2I�e �R2�k�H�	v���)0B�p�A*���¥=���t<��P��iF,�,���2kA�\&-Ծ>� ���Q�z>���z��|�>Z��V]�^3�o�1NQ�p!@b�
c�B�+"�P4M��j$�l�k�D$�0�̈��Ǣc�0���D���R�	y�DILVV4�Qӽ�)yC��K-�I�z[���^|�������g��{G�F����$	I=�"Y:uf����8͔)Í��	�Z�!�]�TiE �*�	,,ҧ#*ɵ ��(��w¸~y�~�O�w�8�|�5��n!w�>ٿ�?o�^�?�RU	1[�Ǐ-�ٌ�M,�QA 4h�-4)���q�(l�=~�}>�f4zr��%
�_HqLu�x����1�o�d)<|w�|����p���lk%�m~�����w� G;����_4�Mu���	�BH@$#fZ�d �V���>���Z�V�\۔G��7JH�bH�MR �n�G�g��TU>_��~e}��}���G�����'��mu�����/�G����O�� ���כ�B�(�RE	�]k��ҪE5�s�����.���5p��ڧ��:%�b���Q�lgnV�OQ�S����\��UgU��6tf%>g�a5x=ݺ!p�Y1���f��J��̪��݋�9�͌�}.'_Eƛ��宿+�xTMí����3���Xa����jf��҈T���	{��까G~��3i,Ȭ�V�W�e��{��hݳ��bs���V	L���7���\v����"��r��J\M-\}>�`{~����HV���4t��梳1da�dܹ2��T��u�u��H�y�p6/0f��ЫDg�vƿ8H[\h\��b�	GG���G��S�2�!�]V]��h��2D�mU��yS;�c�x3�VuvHۆ(��V�G5Чe��̰���5Z�vcs"S��8c���{��\uI�O`cp���|�Te�o�1�O]��K6���U��ѝ�;�v�:n�8���o���v!�dHz!VW�����XfbtF�_n�_<�q}��v>������n�;��,{�i�L�q��IC��4��7
:���V�l,��wX�6UM�J'���]7����d�L��*m2܈Ч8�G�N}kڨ���:$���#���ҷ�uڊ\�Z��d�}L���j�[L8�n�H���@����:�.�ZO0쎼�͜;/K��3�7%9í����֡�p0.![v�V�f��b%vǕ�����o� ?K"� �K��O���K.�[�a��\�M���9�s���.7��+}M�|����N�?Y�=�g|[���T���O���P�E?�g�}{�W����om񌸙
�B~�,٥�*졏�= g��e�CeH�ބ(l���g�)���^���nt�'+�|�uS 7Z��ɱ�-�G>�c��+��/&���$,0�U��Ψ��(~P"����}��(�����uw$"Į�p  􈪜;��j�cȔ��Y�z�*;�:���WN���	Ƭ^��:WnǮ���Ƕ��ݡ`�m��J8��O2��q��:D}��(�j��Z�T��I�|_M��S�	��<�M3�k;���	�!�ƶ-Y%C�n��j���!��/=�n(������0%R�L�o�J�<�=A��	�`���Ҁ?6(O̴�����I
%3i�oQF��h-�y��JL�4��/�iv��\��;���*������%9�S��]��e���z��-��W� c�����`��Vu�V��Ԯ��w���|&��C�Kpfn�u�jY0jK0�u/�Ҿ��7g�$������9ԋ���DRx�sWg�E�n�`�\�nR��;�$�d���> �~�>��e�f��<�w7�(���b �>��څ/�D`1�ʢ��u�g��:�PPX��8��ދ��� v�?p��D��FN>�}9��ds��F(uI&,��I�9C�'���AqIO��v��E\�g���nj�9tky�<p3-hC�xoҞ�f�`,�)�f9߬a	S�W;(<��7u[/6to�:�.U��VUi8�u�G.T��(��/��q.�<��T�8`��s��FY�\,��ˡ�3E�z�$�Ҫ��YQ�J�~f��>U��f^|��_<�N�7y���kvTb�8#9���D�H >L��xv��,��ȕ��]��\��\���h��1u<E�D`�XK�7��t���)}|��l�=�as	�R��Y)M�D�nŭ��z��d���Í�Ȳc���&��迲�h�&���e6�H)Hr�^�"��߇��\�ϰ,��^�6f�TVq��
��\ �n��<v���1IO�}��y$����� P�r��o���&3����%s�h�İ�pk���V\ݡdd�{�ޗ9�eNu� r��$�� {NA$#�%͜���4���+a��@(�0Ł��������K��RU((���ĐEm�W����v2f�P	PqR�'��rD�6�)�u>��h�nP�eεd���bϝZ�aF�C��D�0��!E��Z��^"���Ml���ї�H&P��{��kG�^�!�A�d�����D�(!�aI	4��L�����yD���$]P~����3�q	���U��x̖��Ǎ
4U��00��y"c���)��*�]�z��#���0Հ�Z�Za���Ԙa��f�GBW!Nm㯔&�UqJ\���;��Q����z�Rg]���I�{N����Z�]��-t)��{��u��@�)����4���N�v/��ޢ�Y���Ζy�s���zxfz\�︇�u��s �\�)ݣ)��������G�;�t�*��lN�eL�rL��J�:<�t=S��;�a�%��rȸ+�:%�0x.k<P?�Lf�����3��d���	�WГ�5f�ܹ��NU>~�n�8)!��d�uϛ��'@��F�ڠr�r|"!z�_�LhQ�*>�mg)e�����{�7���l��[z���� =���>7�p#���+�z��?�I��>_��?G�	�������8������-ړ\uHم?cx_~����!��l<c����4�a�G���	<������I�����0���#*$�����'T���h{|S�f�n�����|Z�����k�zA)L�O�챮��L�k�TK�i/�����a�*,D��a
�$��9%A/�L�i�z�&����B��?C����[���=�޷mw��,�����v�XR�cE��	�E<F���m��ahY���h,3�8�j��7G��wH�<x�.�&�5��Jp8JF!�@�Z!�X�.�~r޲X��$'����vg�\�n#>{A=�|ԗ�oZC>��z�o!��.�y����1/���u��S�a��[��->U��k�gL����zZr���C�^��P���G{)����l����Q��D������o�Xћ��I��ϿivJ�E$㦓��R��a�(誰��-�6���H&�������/��Q��=;�h���<�,�gï��Gk�>7�j�=&�i����D��鵽1������=b��G�4��mu�k����e���B����Q�Q]�"jUqFBȂ�  ����4ch��X�0B�U��o��y�c�q��W�:����y�ӣ������z�'v�_/�����;Ok�2� ��y�C
�d/.���tW�2�wce0FJhXBf	 ���M6�!�Z޵��D��R"���x	�����m9~m�XO��~���_�|r1O������=���?����a��u߆������7������b6�����i�O�P�cc��.��&H����3 �====���.���<C��Ľ�/TM���r�ۋ�˧
�b�!a��l��!���Cw=���J��I�}���&��ì��@�p��&���"f�iG��W��N��tQ��b� =��� � � @�=7g!�mK9V�0�u�Կ�C,ɰ����W8O��83~�CF	��/ˠ�4��qزD!�Z] z�H�Lb�+
U�M.��7��٬��J+,��M��](A��4��+�Z����9�ت��S�g�xZ.0�����ҙ+f흼��*����sXt�h[s��LvKo����eƇ�,S��KBuoiZM}�5�uD�9¯A��D�y�\V��!�1�ۄ\�:9F !�=1x`#��-7�Kn"�e&˕�o�2�?Kz���b�1�(Ч�e"��qD�WS�2*:���7Ҫq�L���sS8)�l�wI����!���Y����i8X��bj��wh����M�f=PD1-�by��:T�ur���͕<(Q�"���#�B�8�#��\İ���z6u���m����ma}<��^��ǔm�]t�OA�+[�/tGr�բ���8Ɛ�5�M�rP*eC�����[:��H���@�����SfpK��[F��Pr�8�rA/H���b�g:J&d�%���5O��{��?�`���}�EEp�8�g�*���>�l�,���RN�}q�8�)'�<Mbr��X:���5'X}HC�6���.8��f;?4�sV���ʓ��+cQX�X#4y��Nxԙ��#�z�A<`JD�<��Zԓ�;br�tX�׬T�6��bC=8u��K�k�Ea;l<�S��U�+/U(I6:�y��e�t��C��^�����$�#Y�-�'�'�t3��S���dɡ��y���W��:�[�S��˴�a�
�\(
gd	���v��0�8g��Cn��n�fVl�[MD��֦��]q���Gv/j��,�I�:%�R�τ������u�\�f>�����LERȴ3uR�-�8�����̼���X'a�g�px���.G���yi	�K�H'M�.掫tź�����AU{��!,T.�����U\�)�vMk���_o��)�&P#��m��J
�8���)����S]5
-@��*����+���k62�3�탄蔼�-�M߃Q)��A��b�ۀ��l�!N�ln�ͥX�8&:��y苽Z�2,�9Hη�_/��r�dg^���z�A9r�Ӈ��Q-8�0�rC�g@�'�Y<\��P(p�F���1Mw��L�1��7�#<Т����!لK�)��3͆P��B#s���|~�5�������0���!��H�o�&N&����L뼍���=j�f2�	sԤ��Өp�N����-�V�&�Ȯ=�+@�u4����U�2�����8��@(	������a��hv6^�J���A)�1)#�\7Dz��8��gBFP� P�@a�eNGLt9�+�k��&��T"���9 Ei�1�w-_�pO^Ƌˆ
+���"m.^r�Ԩ��k��KX>�^�v-�JD��\�nnv�r�V�wDp�m;��� �D#o�r��J9��N�Ƌ��P#�;Q�\l�fcZ�B34xMʼ:n,��1��V����V��%��)/?������S����b�|��[y蹢��|?��?��>���,oZ�A�pb����"*��9 ��A���1}������g�V�����X���v������?�����E����w�!���'T�}=��|{�רp��:����
q鯽ϓ�FU�{IG������>��w���緧WK�|�|wA�:۟G􏐃���+�o��ޞvꀌ�{Ҿ(��#���^�<�v���}ny�=��Wܷ���G����p�ǭ{�氈ϟ]���i���"�lVP�����=�#_�Z�e�����	�k�ٗ���}������뿌�����a�m�zv~�l�sνk��C׷�k	����ҭ�U�qis�_����n��qM�c;�-�����XfE��{��ӟ`��z'����N�7Mc�X�`M5|�Yu��tn�u�7��p�K���6��}=%�B�����v�W��w�N��8��"��� ��tn�{��aNa^�~}�li�>�����m�Ɠ��7�\���Z*�t��>+��߈�~��<�(R�����d��m�F&�(�J����Tb��d*I ���۵����U�7��q���������os����_�8o�Y6*�ܐ����?��_�5�VzG���b �#��]+m�::j&zPw&i]�v���иbЌ�	�	[��X;������NVɜ��-N�܏k�iD	���{�{E�b�@�
���fv�a�������S��eFs�0]k���g'����mG�]IS�ەE�y�!�(H�dKkE�Qc���)4
��f�5��*=/l]*냽sK��j.	QHI(^J��UVLP[њ�7IgG�L�,^aQY+9��V�$ڲY@��qq5��9kQS�b`�����Vo�L�Q鳊�N#�'z'3�d���O�TD�AEL��t(9���j`Zw�9�-,|�Ț��j�_]�X�Û0����Em�F���\�>���zJ�p9·�P��U�[KaF
�p�"2���nf(ə�퀧͝�w��u������i�Ul9��0�;6M��ui�q'�\h[�)��������l؅�,�#'kPΎ'�J��m��]��C���`��Ԟ�OnF��f������LP�t�]5�yz	�f�����ش��Bֻzn��Dmb�'P��<FX��9P��7��n'~Qڞ����"�;�cR6�U���Lnɋ�V�S���ؾV�A�c��I���E��5i:��8��8\�]�"	�;�*g'�1�`��t��a��8���G�g�8ߦ�E�Oe��\j��L�eius��F�fc�=zӉ��9@����}���I�y�,��nv�) �VFU�p64O2S���y�^�;{w�0hh��Q3��+�깦f2��ˉ��͹��̫ýq�o'&6�jK�;9=���;�d��c�/z�d��n�
Q�Ni��Vy�*sY=\�ـ���s����aTǚo^P�]H�Z��hOU��OG&c�GQ-�:"y�Wr(V�G�f�%ZrM��X��vNt�|���X�9�uU��|�d٠�Ş|"���y�oJ�b�u��nຊ@�n7�(0��D��1�Y�'�;�Mm����3����/�y;����*�e��9����1�nE�}�>�<�<��./n"n��\sz�{�Tn�f:k$�P��=��Pюf�~u$��B:B{����)�9�}c�a����I�z�w(Z��Pl���W�bNM��YO�,��d^�83jr$ƽ��V�����v�Q����Ʌ�{���T>t&:}��.��ڈ�Km�g=DE��B¦����w;�'�ܥ�J�I��%�s��YdtcGiڎ�Bp0M��/��F��F`���!n�e�U`�
�d[t�d�������V��G'ф<jD��
��]fT�;���Qp�28�v���gM��H�y��uX�p#K����Tt��r��6��X}�%b,�P���"�VcYyV�6��Ѩ�YU5A�3��K�v�G�(r��G9m�L׆Z��J2�M��S���zbF�8̪��Ӫd�t��E̬��Xdu��}s�&+�sja�޻���LPxD\����b�n���5W�[���9:���&o�<��!���ۧ�8N��b�I<�U�%�ۚ}i��n��ޱ�\Yٹ}k#�r�0S�;LA!,�՚�_K��ܺ7��v���{�z�|nIu�ih�x+i�jfk=�W>�E�Pb!+�豵9�&5�tSnk���^EuṢ͙+Ą<���	,�˄��/*f��
�ͻf��vʡ���R��/;N��'{۫N�.`ȨDY�������q���F�-}7�|�tvq��9=R|�xQX��a����b�������ڡ�����B��$��M������y:T�4��ՙ�;ż��w7٤�)�/M�)���zFZ�AT��LI�r��]K�flu۩
���l��oP�ĩEi\fF�*�ʼ'��<ghԌ&*�S��Q<)s���1��-٧ۙ]��fT�sN�'{Xao%�f;ѝ�U_m^rY��T���eFm%{9����ֻz��p&j.��u�o��{�F�mGfP�K+n�<����+.�+q�`����"y�ޥ����7��"籘�R�ٶ�\Iu�u�NR3jr9Y�Ǫ^N:��W2ws�찢-���C63�BTJ[Fs���fI��QkM��Ι�&�ȁ��{y�먦�wR�R��$<3��Odh��`7ri����4�Fb�;�H�!L&U37��ul8�wGiކ�Mq�'�h�ի�"b30M�
��ᦚ�S��'���ynoP��~`��!3g9R1vBUZ��djsw��C]ys�E�n���l��[+�3���T�'�B��w�J���4k�#Y���U�&:�GleNn��iU�����x��*8���:�ma�������Ԑn��*8�D��{��:�̚���{�.v;�Ꚕ)�4r3ti3!Q��Y�r���q���<-��VMQ��다y]���lxr���aF�(x�g7���WDm�	RqҞ��w��"��XE��3�!H�s�nM��-�L�}�1%��·����DN'Q����M�N��8�-�P�m`h)���&4���ޭ˼{�
��t�щ��[Q7xO�qx�˹QOjFF�^s1}9�/l��UĝU\�F��#�r.���N����b�"�謌݁OF؝X-�r*���U<x��H�V�p<zn`QD�w��(�Ѷ�V���%�vs	�*#6�\����^C��;#/���Q�ζ{����O("#ȻvNpק\`X��S��sR�h�����wZ�+��k�>{qr{��.]�7����9rE�f���[�ՍMĂ�W׬�z�tޅ,�Ğ1��Uf��Ag�k�tD�F�E��!wL�-�Ɛ�EFA�:b��ȡ@��m�'�m���i4x�S<�%�g5]c�+P"U��Ħ�*f��fy����oa��R�&�
#��XHp�.$��zm�m
]f�Y��o�R[<~�����y4z=�Z{�b
�ո*�kK{L�;�)Q7I�1UW��#l帎�(��gVɽQHl�����1�2��l��s��jg&�uM�7���#c���7�ksn�m�]y��>���萱��%@����)�s�A҂�ROe]�c�`�@�c`\o�>Ȼ��N>��&�]�8�߶n�����(�!T���T�:�j&ghX��t��vc���p5
�dA�� �"�o����ìN7�so�|����yq���5A��z���&oPi��3;y���0�����U-�[;��M(P��q�YsY�fQ�2v��h��7+��D��[��T,���ЫQ҄no`�%���!��ҧ��V1E
�^O@|�p�s�H����n,�dD�֪�NM-�G7X117�vn������-=T$���뭈{���sjq��1�;���uM��\o6î��=ήw2�b�D�[�vI'����Du]1�#�vQS5�e�0Vo�;����www:sWoIڛg�Ell.�3m�tt���ݡ�y�XK��j0�ս�Z�!��e������	-}{�b����Φ��v����U7]�x��gr������d�\�`��7�ivqVލ݅"вA���	�v����ꩱ��@�j��r��V��{�Zț2��,���YCg*7FKp�N�����K$ĭ�[��xy������yN�nt��ꖤX&�rJ�{��tc��x�&��A��ߖ_K�ԱWm�Z	ne���6���J�bK�y樏Z�I��Zk���o���9I�q�������k&6#�u��{�nV�y�C�D����%d��繕�M�=U�j:�� ��7U][S>M95`)���7�.ٻ��{�'Hq�3Mm�j�" �\���9�a�BA�U۷7�gyT���ݖ��|M{�JX�욫�'�RB��D]�=M��Q=}�Pѵu�&,疠cvf-�j���ݎ���}�Q0�c�l��D�P��[Aa�I��$��J�u�1���q� T�����!mU��*�q�];I�̫��ݗil�*2�Qu��{W�Ur. �nB�܍����c��%gaL�*-�����f.��`���uM�� �9MD�W)3EOq@�F�a����I��5�4�
�9���@uGB��8�|�P���&�Y6���F��w
m���q0y��k�\kih\n�̖����o^>����c���zV�p��wU,�Tf
���x�9��r�ź��v
���ٍzN�֯`9Fƪ=����DFe���Ry��T�Wq;�*ؘ��,9�2�i��2�Ϛ�:��l��2v�WN�Vy4�7��ɊD�#Y^9؜@ȥ�g�H���0e����j{�y�qdW�j.�cXG���[x���s9�싙������O����ǹ�P�f�|�J^��,jQ����.5���o�(j�*��ʪR�WmfE\����F�;��^��Q�8��~�����qq����X�LB��C�l��݋��&dҞ�K�Z�S�d�Y�o������9j�*�P&�������m9������wn���Yܩ(0Ev�v,��Qa��gQ1]L$�e�x�:�u�Z�]SX&�Ic�^d�TU��]�U���~�?UG�\CI��O*�О^��7"�����9n��nu]�C\*������ad�7Z��Lq&�s,����5�Gm[��t�u�Ø<���;��T�|��% ����c�.Y�˝�l�Op�[�S4ɼ�
�K�N��Ұhd�m!�D���4:#g![Y����٬U��ٜ3S�w0�f�5�+TjI�#Kz�������0^L��3�hQs��eq���"&i�b��G�J���F���������0����E=�V4%�<�w����'o/�ciN�-̾uW5���J�v )�f��ˈ����]t6k��'7��t��^>=�����^���[�)���V\�1ǃ�5O.6:v�$ُw�;�����;9p6k,�p��3�&ΐ��q���O;�ђ
f��T�1Q�ơ+�%v����Fp�]|����U^L��Alb��̾�OZ+8l]-�<�����U.ir��vr+s_�U�h�3l�r���N�Y��V�f,�ߝ9Ix�tX�8�1ұ��lf���]Q]B�`Q]qS�S�q����cI�T틚�����6�CC{����U2��VLIs75��Ŧk)�Q���e�]����r�f��7Tq.fghn��X:��#p�9�J]�eN�i��ud�wK�T��t�3$J�9����;d-ŷ�*�`��B�kz��Gi�����P/��o�w�aT{��c̒����ʼ����b؎�rdZ��y�ه�r��'�Wb����"1���&NU]B���X��hg`"72�p��k#����3��6�?:fS)��j�N���Q��.�{1X=���$���g1_�w�bx�5./]��F�B�/_d�f��(T��r�_T�m�۝�'��v:���� C���E�OL�������U�V����Jp��wE�n��%b\���;�Λ�X����dÅ�5��ؾ�3-e�]`3ѷ�����%pu�8{3ڊ�p�B���߭j�9y0�K�$���vx����j����ˑn�n��"'A�{g>ٗ���H?q_��L�܉pwG<!A����@����9亽�N�8���VX���Swv�8Ɏ؜Ȋ��u.N��1\�g�N]��S�Uu��I܍�C ��Dm�	�y$FE�ӹKzZj�\Y�7��a�䣝��o����kJ4���m�h{V"w�ނz��{{7����cz��\�(:lLc�(�!֩��#D���`���϶q�}�8���5��p�.2.������(h��;��)��F2�K������d-�(@Fkyu�6�Zޓ/C�)]�ꇪx�qc�"'��0�)�Qv�Hr�2���e���W9�������Cef>���p)K'עa��$\��3��3��;f�]���'F��,���
���J3�yTP��t:-��85ub���l;��iַ����z�TS��St;Tbw�J����YT����J۞B�c4��q�M�N�%��wI��m��x��T��,k�Y�g�b64D,�Q槕���l/qtVv�p��Y^�z�f׾�X}۵[]�q�{��:�_l�\P�*�bSGw0���8�6c�6�ɮj�3���m	yu; �na�Xl��ر�����d�6�)�GTB��U�	�Q[㡓�V)�@�UO\��1F8�� ��R�97���d�LRL�u{o.;�k5^�׾��B=�<{D���˒��3�*�L�ݦ�M��]Y!�̜(藼0Hǂ2#gA�dU]m�fK7�Nؕ�UX��h��,`A��{7���8v�*���F��[uG�$s��gP��X6%@�mI�ŵ����[�g�ۇeѻ$&S�-��b�i�V�eM@7=ɼ��W6�yمt�f)$�UV(��rp���uڌEV0ﳱj�RN��.|z���ٹ�O+g)��F7���w����曬��J�_l v��Qٔ�F�{�|cvqP,�;D��,]g#՗JN�mU�S��C�\(ͫ':�'ƌPj��z�)Ѧ�Wkn)�[�rѵr,�F�J�ri�<(<�Yc�ch�[����ݞ���_:yHdf��gkQ�=��d���ݩ�4��R���z�_`����f��lQ������$�k�aO{�������ZY�N�s�iF3Jy�b�ט/�5ra\��
����gd��q���V�e�8�tF�}O��ٺ��EdHTO]ϔ�7�s���f+żf66:�1�#T��ʻ���j��W�ҥk�M5Kvd\˱�N3�;Z^Ou�Jo��lL͝���n�7 �nV�]��������w6�ꖊ�1��ص�MR�'k���u�W��	��}p�vi#S;k������Hλ�%30�f�H�9�J=�<�f�����79�D	�8f��gL[��5�D�Z�=�jw�R�ğ+,hԴEĭ�f
Q2���+'DMƨ�̽�tpXw��&4�]ʍwz��n&��\�ǔZtuq:�[X�9(O2'�Rɪ*�E�^!s⺱$��}g�S�ҶAܪ��|�\����g��잁���.�v�Nb[�WweVps,�z=�et�Cm�˳�H�q�D�����Q9�f��O7�*b�D��/��E���r��R�w���`��jM�����;��8��\d&0�T&^-�0B�Q�����Ⱦ\P�vȨ�9�f���\t��owp8#7yB�u8����b�f�����:��ٷ�;MwR��G���<��p+;7V7/�(�J�/t�{����oÁ5�{H�Js6 k�Y�l>�}ݹ��G��TJ��v��S��)���5Eq�R�zJ�.5�_]�i�3�U}�Ή2���+�-q�Ԙ����؎�p��[z`k1h�0�@���]:����<i�i�_���9�Ĉu�f�k7Q���;���y���t�yFzv����s�7Q�t��Rdt�8��*뒃J����e����EfQH��α5[1���v�4��;%�L�h5Aa��W���VBٓr�V��B�e��Ds7�iSSb�:�_[�B�'�]Gp�����fb�E&�IZ^��^���:bjM�׬my�r�o�U�×�n���
ɩe^�M��P���3y���[E9;�5_n��;��}��m�&�O�3�N��l��� ��jMS��B�5s�4֊P�l�3f��G;�+��rj�9��ˍ��t1Z"��_n�4b�o��"� ﹶ^�;@�|z"�'�)v(f�{�3Q��Uf�1
َ�"��ǋ���-�l�Cw�g�q���ΊU�7:�Vu�͋��*�w�RZwtZ����k��m����`鱕w<mM𹭩��Sސ�y�q�^)���o�B�p�S �D�ؘ�N֛�0]eż���:U)�����7��=�7=钅*O�'���9Z��9oh�����T�Qp�XY-�ۘ�Ng9���&��qSyO��`��]1_iۻ!	���2�.j$�f��\qs�|��X��{r-B	+���%�@�U'E��J����1l*�G��2���-ٝݫ��2ƺ��xaS��ͼ��"�j�`��V�gn^r����EӮ�Q]��F�m�2���U���u��]��.,h�]��4���E��lD�={�B��f����lȣ�D�ᢴ����㷉���i�,a�p�!�O6�e1�$����l�*7�`�N�������3����Pvd�u�u�/:(�+h=�}�	M���gsjgtl�����+l<�y�/W�b�����ՙY#z&�h��bⱽ���z�񉄶��4đy�A@ᜁ�v��Ggޚ����m.؜Fy�L�rk�zt�[�]�~ڂ\B�HJ��N_O��C�UW�q��"��[�W-��IG�³i
����D8���(�sAZ�����u�6���Π��y.ըu�OT�Ko�C.�熺*�VM]�J��.�w��a'�y�38ƹ����w8�7S\��fv7�����Ja|�݌문8�;�Ңb f�y����'/�:n��5��=���ek�ћ�2/g/"�Lv���r��v����ی+fk��l�Hxz�+F�*��
c!��K*��	r���.���|:��Y[*�-�}�m�{=�N]H�3�2�P�.�^S�{�9���`3�N�wN*��5�8�q�g8��0��oVA]3�SW��(w��U�n�6��bj�{t��&��L��P���:4� \7�Y��!�����Tͪ��=�{�s�f�OEFh�8,a����ND�݀��K���}9�C.ᨖ���nVԲʢ�E;vv�I�}�ugn�p�ښ"���3�0jQQ�;�\:='��_W���a��O���S~����)��^��*� �wo�:��Z7-�C	�E�������]�P;N�҆�\E�P��Ґė%/7�as}�>N��K�m�-;�Y:{c�غͼ��V1w1�p��KR���q�5-�*lq��r��1�m7�͞��3��[g2�y�8�O@�t �D]�1Ӝ��fv�Q�3��p_�w�W�~𘲄6n��W�)��[�}r�t쩋Vy#����3s�;�4�ź3]�7�Fܿg͜ѣ��~�A��v�k�{�:�*�d�(<�AҙZ(�m��k��dm�9�:͔1m�9¿LAy������ET&jdҎ���q���N��Q�̇-;2,�'n��nF���=ׯ�W==��=��[n��0R���>B��p�z��rva�v�u(�NÝ�p:�U_[���4D�y��B�����\���=2��,�鋋A�Wy��ҹ�	��Ei�[��;ԯ�3r��j�[�f<�ۏ4Ml�J�95��Kzݾ=v��؄!͢�v�ۖ��Qs�L<"�0�]l�Eͩ�Z����M�Y}�X"��d�aj_*�DΨ�����6'���ut��˭����f�ԭpG3Av�F�WR�V�����F��J�Cт2{��WT��&u��H�6���boq�xh��B0r��z�[Il%=�.77,�WE�."�;\ts�u���y�����1e�i����^��Ε�Kޭ�o,Jiom��YZ8l<�=z�;3w�8ك�z�Oj9u��d�����W�;z=N�����lc3{]��m��v0=���];�u�{R,����l\��)d匞��U�0(\M���^���V�lN_Wl���������6�39;&�\乫�ivs���ǌ���*N���3.�3Mo"vBެX��p��y5�VTe�}��'�j=�{��Q}�}��.5e��uf�c��=!)�W={.�EG�ʨ���Z�n��mgQ�9Phj)f��j��.7�kg���	ueɾ��{�=§�����{�x�D���g*D�lU<�tv!;\�O�(����''�9��:��wE��Y������{��7bs&��c�o�+���Bf2���z�:�ʬq�������A����뙳��W+���*��l�l�j�S�" #*�"HȰ��T�c[W-V�J�pۛs\��k�鵒�wG6�X�RM��sb钭�K�r�\��5;:K����D-�\̃KVld����\ۺ�k����lEp����H�]w0���w.�u�\��M��N�n�����nc�k�6�n"M i��b���54���\�4AL�
e����wG"��%�,X�� wG(,�v�b!+���P)M��f�lce.��dەԂ�cC��hB�;��d�͹��-��wr�Ŋ�7uһ�wh���)���TknX��r��IY��Rb�خZ��1l�ۑ��H�uu1gq˝ݺ[���ȫ��r�v�-�����5®F�b��m;��1��r7(�v��#q����'v�N��WH�v�Q�θ�m����t��,b�].�ۛ��M�nG�>��-d�Z�Օ�	 �G�6\W��'�s����t��}ur<�����,�!\����{�m����/iBo|��_z�ޯ��q({�XyT=�'��=�+�B�}�A�x== �o���6�BPS�
<ߧ����Uω�C�E!B�����*!��m��/sʐ�j%���Jo���6�BF�%�HgrGƝ��I�ܭ�'�kePd����s�B��i^15��G���!]�//�J�zz���\����7[�1bY���ܭ�Hh}z��cx�*r��b�Kì���<���E�S��*���\v6�'�"f�oX�$�Ƌ<Uܻ����8�W�YDN��AN�X|V�F2�1P��))�ZC�9��v�=����x�G�L7nS��p^�R�w��[4o<�D4̂�;oR�Cy�cL�7�"�ɋ[�F�i�]s�K<!3*1����1��4�G0xN��2�6��d
��M��Տ3�<�\���bmZ�i]�c=�˵���h"�:�!�u܎}�����Q�<� �d1<A[Gv��V=�\ƺ2e�xs,r��h��_X��m{��E]��*$[!E-<�&��;J/�u�r���1}$��D���ͱ���n�/��-� i\|��ij9%?:���~/x�&�*660���4���\�:�� �b܃9��y���o:z�o8|Å��Y~8�T����:2�z*-mǃ�5vq �i����̢>��3��wm�If�c��V��d#���e��5e�N�����]���|�o�R	�K��whT�-U�.�(����(]r��5�T�7�{�F�^uF+�o9��*�/"A#�xb���bN��
�������d5�5���m \�"��H�EG�34�+M�0��:��)y��KG��f���C�2ݎ7`<3,��p����t�I�){I}"��J'-��~=����� N��^��/2�Gj���-�%!���܉ֲ�^�[��uc��a���.y���z���oXӚ��ϟ,��I�~��8��"		���שB�ߏt�{.}yh���2���_U������.�Ľ��:��� {�3N>O���6�E�׼�@�u���D�W�ڙ�d��9Z�������=Vx�-���x�\e��S� ZK���v!h0+��Ӆ�Ѷ!d���u�a�N�~�p�:�0�ǥ'�*�kʴ!���]Ţ;��~��&�Le��Ҽ� �ݪ��q)���������K�C䫧��0�U�u��<̯�ig<Z��A��5L�؋�p_�
�Fy���d�rf��	$��#�A4��|���d����:�o4��B�=\��H?F�ٮյԗ����ᮏe��Q~{?�8�D�yٗ�ܢ��*0VOH���h�bF�б-U'�h�!�x�C֣LsNL�)��5��;=��깎�;���d��u�a�앾#w"��j�i���F�* 8��in>&�j�	��]�$���@�rN���c���?%�s��D!���sT^��Y�"�J%Ķ`G��x�x�*ԁ2�F��b���^Y��쉧T�j��Y�c���E���Ɨi��G.����N�|�9��R���Pd��k���;���B���#ܺ<K	4�'�n�q���NBY"��	���N�1�nOy���	=��F`g�"	Rb���OJ�&��I����p�����p������u�	�ԭ!��
�71	�@�3ᛯ�*��vl�,���z�����������������~�B��� R�� �
8b��͗�#���H濭��h�~���Mk���~.���9xj��S��s���/�۪W���(�/��e'-y���D�6ߌ������+�idy���g�R���/�̲:'�����8�Y�Zx��x�T+�N_ޭ8w�7�^����ʯ�/Z3�wnݺ:W���k2�uޔ����/<?����Wi7{4;��m��3�����{���]�C�����������7��:���i�n6�o?Ysy�}���m{i��k@��%��ɿ�W�z/�kq��3Z�ͼӴ{����xI��k(,#�H��V���hm���]�>to_3�x�HF�$<e���zR���6�����t�<�"�g����E��!R�)�����^(�� z�	 ��#"2+HKEN���?��?2y�/������W!���_��?��rw|���yl��W���ˎۑ|f�Po" ��܃b(�NC��|��||g��9.��Z_��k����;�;�����=o� �l���_.��۾�.|R{�s��{C=���d��ϰ���2B/ѼIƋ��~>������&S���'�a"���V5��[����-�0̔�-t��>?/��v����������9��LQ^�t�!e]��F~�����K�[� ���g�WMԠڄ��#��w��~�z���>9��"F�g�35�J�����S��ۑ^}@�ug�{bڲ���z q��'1��<���4�%�ߔ��-�l#��e^m��;LpG�p���i$�Fn�8�H��@�~edB��S:�����ret�1�Mӷ[2
�9l���霈�F��,:�\��y����΀�?�Lg/�����	U�.�>^��1��K��4�V��� 0'��@�0�Tx0S��L���DB6n��röF���0�T�HS�@���ˊ_T	�+r���Q$���P���u
�Ve�U~�!.���V'����%S����!�(�P��y�Χqr�Ŕ�U}I��2��@.�88�>��|�_H��q�Mt]����oM���F}O�7#�Jn��������Q	��ⱓ��)�k�V~Ϸz��%|�1U0l�P+��\�X/�#J^M�k&yf������xZ{ͦ�ٳ��Z���t�ʦ.��Y>#nJJ�N���ܳ�gH1���ʲݵW����T/ ���N�{���^���8���d�s�0��Ѓ��l3�L�~X�ڜ�
�O�g�D�G�A��)�?99�b���l�k���������
q1\�;�d�J�t<̷7P����-�g�O1�n�^z�,�a�]����MX+�j7It�#���X gNd���Ϝx���s�&q�{{cܞd9ɪ�VLeӣ=Ϡ�<r�3G���I�����N���w�1~�󧆉��:�/�s�ͪ@�RH� ��ݢ�4�C�G�}2�
4��'���:�Z;o�w�$�ڣ�p
��W��`.L�״�Ͷ�q�-�����w��s@�EVi9#�p����l�
-{�^�Lw^��!�S����s�&��9�'�b�U���z����E�[Ͷh�.X��/�om���Rrq����Ø��9v�#�i/rL�g�vdu�1����쭞T�BH�)sC���~�V��p.e\��w� ���Zwl��]9�U�z�����Ħ�nQ���QR�9T����E�<Z��0��w����e��3�$��E8��d'��=�л�!#SWs;�����Q�����(��r��=&���=؍j)�DS�g%
Z7��^�;Ng�+/���2��c&�;����Oy��+`Z������;<��9C�x�M����}�N�9�T\ޏo����Y��F��qr�8a��\*��<�ayz��6Њ�
#[�'�N@��{<�7u�T<��i�_W=Q���� ����e|`g�f�o)8��P���j��T��%�-�;��R�(��t����������=q�y�;綔�����>IEX��sc�G�^�'��:Y����b�����9���iuF�ZhMV���9t��|\�e�DV:�/A���S��V�ؓH�ǁ�40��hc }��e�i�u�bq^�����8t�z��O(�Q�^�d�`����fײ�[�͏�	������l��D���H���c��  ��}P�9ņ.b�!�_����,�T/���v�}s�x~�@H2��[ݡ��g���!�ծ?rῨ���2���4�Y7�\.��8����J@龺EﭴM�f�om�F�S�,���uXTBO�
r�i�p9�w/Mm>7����:Т�st�C�b#%���A9�
L�s{�Vק�)	�W�//ۮt�ϝ�\C\u4cRΜR5G�!Y>k4x^tE�����w�Mٱ��~��FIU�ţN��NIk'�i�W��H�0�i�:�\l����F��Ny�l�s%��-�\/,�:���h��KS�¿��M�{'[�r�y���gt�w�Sh�$�:���x�Z3Nϲ��A3����&t�����ȕ`���il�;��N��$���&�������0 F1A(�50GEj �A�KAQOQ���<Ϲ�۷���'�:�����v����9����r�>��m��M��#m��S��PY �I	!#$�� �����o�m���,x���rnփW����)i>��~c��������Z���|�ZdE�k\mII���'LN��)��mL�'����Q�%b['=!�T]�����k����,�{�Z(}H��"��Ak�c=v���m��/��vh�uՕ����C,��]D�y�Q����K:$�`>�Κ�:�5��Q�j��1~���ih�5�i�kj��z�!a)d��]��j���4)�z���8�4C�,��� �/|��F����}����&nna���Һ` �d3�x�s�Y2*� rb��M]"�'��5���?��v��|����zޓ�u���+��~��k>�����)� �e��
�� R$U��R
A)H�b� �EHd�7�zD2�A�.��V�6ƈ` � �N8B�# �9c��)8�*`�K�Db�4eW�pĉ����R�t���nf6'᯵�O�¯~�I��K	AR��֨.'t�䐓R�n�j��|�A�z]���byo����������(��v�Й�d�0u٠�]嗿Bڽ]U_n�)�����f���Z� �#+5�Z�+����F|�;U-*V�m q!����tP@z?�w�I�Ă�"&��w�2X����������w=7�;O���Q�ײ�=_m��_K�p�_Y��k�-s�����U�ފ��1E*R�DS~�굦������	3O��~}�0v�Ȧ"o���`bU�s��$��_s6J�e\�姵Nw��mE�vE�4K�f��ȫa�WlI��v��;�&(��8�Я���i�J��K�ٚ"�jf?@�f�$�� .i@o�I���x�����������;��]�9?�:�7��~���|�_��O�P6��@��(�6`D����Fl5g�vY�5�3N�+�u��{I�<{{�mm��;�N�λ�U��;��6�B{�'n��+�^�7����%ޭ�<wxݗ���$�~�L�@'�������1�!����]!y����K�a��$&�Q�jũ�ӌ�F�ԚYY��>
k�Ɛ6���n6�U���_��>"���6ƵHR5u-����tJ��s���6�ʥA~�J�rЁzBz\���`�gWa�8U��XZ�tA�߶�nkl�Ϭ|5�D�&Mj��As�"��{��v؈�D"���F����7ڡ�8��G=t(�C~h�1��e����������۶r{�%+}Bn�\Ȫ#�yڱ�7��[-�I8z=��C�1IvIN� �T+
c#L������Qk���[�kX�"��| bT��!��Q!�G��=����K%{�����fc%H"40j�}�Q�l,�tU&E1F"�E��{����K^BKH�©h�/�(�q��:�.�15R�-�0��zI���ˉ6�q�>-GHV�xD�Y�T�<�&�>`���N+��Is�]�ٛC}"Iʾ����or�z��s&!��8�h�ջ�T�u���/,�zV��(i���Z�ѕ�#���EvR�!�� �Φ��Y��5�b�q��8@�؈�Ȑ���I%*�4�(�����ct�F�������|3�oQkɭd��GA�+j1�dZ�d��^w0|Q�*+����������?����������|�8U>$��)AQQ�N݊"��?8�A��x���LA��IU}��$�+N�-�J��\B�.����DK]`��zc��q�Yrt�M��D/��L�U�����(�pD��X.���d��,E�;�V��Si �x*��36Wk���3�i ������=9�w���?�Q��(@b��A��~.&/T&hl��.�*���)�R���z� /�^F{�n�RrU��C1@5d�?	Q�u��u��j�c������DZZ��x$e���g|�^iт^����:O%�)3q�6����""�֣]X�m��(Z"����z"|HE��E���;�;���}rJ*��'�:,��j���	t߱��A�f2��~��֚름^�YqxIe��L�&+K�$X�$$�CCRP2�r�}-+XWB�Ad�+�q���
�r���R�;�Κ�B�Ά���3�.��&��jE�DWM�8��ʮ�ML��bS�p-�;��4d�������DF8��GZgv:A8�����	m�Ț��*ڐ� *_h�Z��kw� RSVU�[5�3����d�ԉ�:
��Eԡ�'LZKG��D�H�0�gs�lD �3*J]-Չc��F�����*ˌ4;�4Bs�4js�_������v��򑶇x< �x/�q�4��=E�z��dD���W��&��a�n��,L��Ќ�"�M~�&1y�XJs��Z�3�đS21͡Y�����񑥀�&.�D�P�|���ͣ���ű�F��w�U#��aPE��P�;����v���X��x��p��5�|�B�T{�kM))�Ғ����t\��r�$ན���i�[$nw!g'���l�ȃNx8+�c�(c�}D^��w!ޮ�ǧ[~��m�h�v���:���S���4�0���1ل`0:M�P-;Z	d���"����HN;�a9 LZb�/��κ>7���E���0!"bn,3,�<^�.���娀|��0^N������$��R�D(4w���$ 
��"�/ ��jv��m^�϶w���V��5��ЏZ�^Pt�t�Q�<�F�n�P����z2GH��5y, ��͌����I��w�����YsI�#�H>�"fϗ�������1�@n��B4�Y��K�@����'�	���ّJg�]Mל���0Ӳ_ �����|���e��bf={���4������ԍ��-9!�ې�K��*���kjLY�/~m�H�X�'����wC�;��˪�WÁE�h�CT��@��b��aY���|X���P��B����^�p�QB⏗Qp�V�NN"�8#8���&(��~RcI	�txzE�4�Xv���iR��.#ٯ_B�W�<���-D=��2y�Cz�׎
&�L�(P�	g���ض�����*�������C��!�C��q����$S�?,�������+3�Q�
���#m�ͨ,L������T�,��D��T��8���{[�UK߬{��mp��X�̳�x?'LW 
`��E޲�u.�ܓz*"/����դ;�G�����W^5�.�[k��P	!���ϖ� L��LϞco�ﶘ���i�TK� \Tb!�k���A4t�^����4S���O�zؤPFP�������h�+'2��28�it(�a!�.t-X!$�b^��;��vѵ7�0���̐ڡ�؉��:G�4������&�I�A�+�F���B�~�˻�vǗ�v�s(I$'�RH1(@NϘ�E�;TODz/l9!��H/W��I���r���ʢ���(�5��0�ET���+�&p8��]�m�FX�]��j�L�X)�s}�j(�$!��xkUG3��~#�z��5�g����/(bP��$6�t�kg��� C�j�!mg+tڥ��'�5��b��6B3;�j:6���ֽ��g��V-�\;A�[��:�`Đ��t�K~�j8|	6�"D.�dnAX�1(�ʊ{=��mASZ�E�s`TB���ԤP�	rv�S{	U+�&#��8X�n1{����[ $nH.�
��`���� �-o��'8��B�!=�n]~_�ވ0UB9U�G^�x��JP<��Z���� ��0.�.&>�F����W)ϙu��;LM�53D��r�9�^I.#(Ե�9� ��+:���Ӷ�.���1�6TjB1�1��4��0z��J����@j�BI#!#C
�f(.�B.e�V��2�g2��J��bn�\K�zzau���0$�W�a��e��;:�C��6R��*P5\Z��%H�t�jB����@�wnP ��
4�D��2.C�H�V��q���ir�	�PU�$%�z�UX�$
�!q!),�G=�{�/2N	��4@��QAqG��EU��BIETxC��oi
��=�QV/ٖ��"���
��TI�NA]�	S�L�$�?��\�Wˇ�����r��xQ�7�@�+.�@��9�4��	Ĥ"fC�s�{�/�xDC
B�.��I�QnP�P�.���A�
��L&��mk��H���n/"�@@UDQ#Z�x�8��f,��TR�# ��r�Q��G4���X���߷��X��<���z򠚊V��52+1B�I��u�_�j��'����U[��A6�zO�7.����`w�J 2YJ#���>"Z�GO�����DM�"�����a(롭��k;:�5<�iF$0�h9�ddleeW3-K5\@�y+��@dh�"O->Z�����>x{�+�c-��^MAڌ�P��(�M�l��xO�"h�J	�GB>��s��?$��D�	�+�Y���v	~��) �R/(�Рm��w�FTG�(�	p(�3�F3��E��@S�8�L���Hb�����*��PT��:qCeb �@�T��g�=h� �(Q'�9�T ��h�z�K~�>&�� ���F��&P6��k��6h�7�[�K�UB	V��E]��+�3f�cJ�o����n�Z���<�ߣ�x��K<ߦ����.G���+�#2WJ�L�J�x%�MQQ�8�R&�˔P@5���L���IJ"A�g-��QN�:k���6
�YR�b��u��I{�ofL�1,Br��R�X�t�(�B�g.��D�PJh�t���¿�[B*�Q˅sH7dY��g�a�w��KH�E�Agٽw9_/?Z�Gx4tz�=
�сX"�n70���5r����	����,)����v�^ȐRa����B�f@�*�t��x�prtq��E'ذS���Z(��`�"5
��Y	T��KjZ�R��\fR	R&��+FD�U�nEĔ *���63yKA�0��_|?�_c�j��?���L�G�ͪ�e��P'�)������ď:&Ď�ꍄ�GfD-�y	ZBP����֝ ���u�Z�)M�Rb`�X.���D[��F���K���˶J�!�0�XT�z���Ó��V�ȕP�%3R���>Pg$�h��A���TUU �@P�VȉK��aL>4Ol���l#�B��|�xL��8%p�0lV�BMo�Y^/��b	8/��^AEG��Ԛ��4�ϭ!��j��թ�*3�$gg����P�����P�zEV	�$_�`	��cCC;��%����	�PE0�-YS����~�Y � �$[�"�	��)�U��#A���k�]��O	��(��}�IF�'�w�=��/�}ݠ��]<^��")�k*�R���@��)�ƭMq��3T�h�*�[��kX	ԑ7�X$���-)h��{�e�B�A���� 4+fb�M��D�0��z�+(4��U-)y����J[Ih���.+�8�嵾(��nS�:�mtRH�I�`R�Q�O7�|N��I�X�TFD%0���M �� ��\�h��e�ib�$�fr*�%�&����@k�$�!J*͑��5lnو��3b�	�ZUH<�+��%I'�#Ri���/[/��Iֹjt�ͶbxŘ9�|@SMt �����\,�e��������3ֽ�w,�n�rykCN�ӿ�q^�EΨ�R��(ָ~ZQ�CgSTm����.x}���r�{���E|,f�bK�!�D@G$dI�j�v�c��K�Rw�-�@h�L]!q4p��Q�L�x�U�}��{^�h����d���A	a�zVr�,���u[�m���l���F�a��+���1��	�¿H(gƏw�D'�T�@H����^���sFW�J�2��<�5%t��t�mY �}D� 1�x�L ����9����.�HJ�b��Gd�����}�d�X��	�˄!��w��"�jo�J4�R��K�F��M���3:�P�H8��Y��i�X6��$<�}�5��]4R�qGDQXv30�("��0LM�9%�A%���vE�o쵰	���
>��Q�8���y!�}���ނ}���y�	~�
�$e1n�0q���т>׵uLbw:^�{ළ�Gb�����J��*�+��Uz��@���$蘡t�rEE:�v�>y�0�(�yD6��(�ii�%ɍ�p�-^��!j�n�x�+�;$D���B��$�+J%J��0`P��K�Z���5��oT�������5NjN=��b�*��i��)���p��宒i5��/k���H_JA�ʮg�
�J�mMyHRE��m��]�4q�ϑ�k#���H VA,/��jwY�d/-J���ϱ��[d@��ļ&��I�6i,��:K�"�I�1$V|��U����ƙm0��.���]
��;Ft�)�|�ݞ��mj���X�A9�1-TR�qs�B������TْօP�D�E�"��0-�ZFU"iP.�U �l�F�K����G��sXG�2�[�g�X�j�"���$����OWhov�%F���H�g�ƙ���H2�V��A�c�'I�A�b{>�PӢ)�WY�H+��m���B�W����
#�-�g�A����c,`��n�����q������lN	`�UՕ�#���Ru����!ZWJ����HPL��� ���i7�l�,�1Qu��	��,���� ��z[��.��g��~�*���8���~�T��d!"�������c��i;��F9%`�N.!�C*�֒������X��1~<�ч�F(�e�#�h��hTq߆���t�>��H�B�"#�əx�%;�a�*���n�\(����)��҄��B���a1	���B���(�xE�BJ+�e9��'Ga(�@�nr��h�"�$Rj' ��C,4m9��J�b(��P5+e��3Q�]Ml��j�D��^�Z�XLW!�H�jY�N5��0���a�| VQ����^���H�{3�0���Ab����,��_j7w|( ���3��Vأ"N�0^�e�ԂZ�5e�E^</������ϛ.��b 	UW&v����׏��}>��0QJ]��Z�aM�3�YM����t�]x�S�Y�6(B$�����kV��":M��:�9�X�I�M��M�����Q�WN�����M��)X>�W���X��	��@h�3���6�p��5;(��A\�g�=�� ׿m�����i]3�D��K
Xr4Ӹ�i�JA���GY�qN����t���zݑ���j����|B�N�݁��>��ֹ1K���7�\4)���� ���h�1C5CK%�E!��&�V�`���J��!��@�F��Qe��J1ж2�0W��Xm�sh1�jl�*lLM�f����F�R�z�.��Am����Ĵ�NϱH݆r�F�7��Ag�b��$��u��b�&�I��,x�'M�t@g;����]�$�	@j��1���@�
�M_V-���G�s�a	����㨉�a&�]����D�-J�@G�Cn:yX�m����MHAFD@���I^&P}3n
�\`ԥ�]q�i(�1�(�4��D�B�"���l[|o��w��A!�^5x(l��M Q"�b�ԉ�����
씃>�w�\$��[��_*߰������0��+��"����ƴ�5��KY-u�#�Dc��9O��Y">"v�ˍ��E�J�t�iT%�	3*�{۶1ZN�J$@��xγfMt�n�*N�jyg�HƲ�Mp67�S���"��gf�![�i{j�A�Y�-�Y�cGj]Z��2��ty�Ĵe��q3����F�3X�0��&��Y�L��<��ظ&����93^�q��I�������5�[c@vL�C��l�ɒ@�D%�O���˧l��i�"�Dl��-��]Sa��d|ix<@'h���U܈|w�+�a]#Ja��u����h4���������W	NtS�����Y\K����&hP��+V��C1K��\W5�^�-u�p�q\C��Y-b�U-G���PG����h(kE�X�}�ؓl����z«bU�T[XV��p��d�nNPժ`��z��TH�~/�Y�Z�C��m�/�-���{����Wﺒ"T$�����H`��L���h4{�=�g;Z�hU$5� �x�C$�{sm~�h�n)Q`�:eH� �Cu�K��v�ŔU�D�e2��d�Y1�4�e�7��(2��F^�	�٥�I)*E�k%3��V�ar�!�*4V\�Z�j���(Q�Q�pN
,�cj�C�U}C�4�w�m����:^H ��5�j�m�"���il�n�\�	�����i�(.��z5^��Y�k�l�\��X��!���U��4�X٭��~��!@�
GO��#��b7u�I���LY�<����]�#��ײYj9΁S�~��5�i�q����F���Z��ʎ.�-�(����4ӭ$ �����7�E�LJPe��ķ���ʰ��sc�k����mY�\�UgX)���~�j���^s������5C�I;AC����aGV� �M�-�ܮ�ɺ��k�>��C5��/dvҫ�x��ќd��J^Z����g,�ģ��ϥ�M�3��
)T֚"Pd��J�hn�]tѱX���b���Du���l�L����b)���%� ��M�
UV8�iY��x�,�E2�k��7�̙��{�j�*/D�9l}l����Ma��- V��@����|͈Dd/:��4�C1�:�r�uRԫaV�-��X��*�x���bBD�B4A� @\]G���Tc������u����0+c�G/�u�v÷��9/���Y�Ai	�����Y+����.w;�Ƽv�A�"	ɩ�
v�����D#�q�'|-qk�$SlL(�	#*E�
�*�Dc_�ORNx�BF1����&r)H�SH���4"�JJ�A�c	��5�"��F�N�$[Aύt�R�Ѓ����LWB����Ԥ�U�3vGO5
R������ņ�����TqD�̮	-9��`Oz;&R�´(�ֱ��1k;&�)�x\G��h�.;&�\�"0Y� �B
���vL�ϭ㋹�Ŕ����O[�a;2*�������ɍ������;o�b�UM��i����`��\l�0[5��τ^nm��q�\I��*-L�s���	�+.w�	0/~�j4���QZh�=�*�x��
�q�gzR�a֐}!!=�����3�n�3�J&^I<�� ����e�L޸ʎ2�M1	�e�յ�:9���]�-,Ė ��9С*�Ӭ뮷�v0��	�vK�9N�*I��M��<\��fG�+�1Q�[���9�1� &{��gk���{�Q���$�BvF|� HJ��`A��_FQ�B+�)��E�DP�ՠ�P�B�	Q(��l>��
Ϝ}��z�<�@s�~,�SB5�z��ء�*	��DD�r^c�,D]X�`�K� 5T��*41���ԜF�0��J��o�qJR-�x�7�no�D�m�B��k��[�s �����R�# �j�!O��q��K�XOe��lEP��c]}m9�uV[%_uu�!x���g�o8�݆Hɂ"f"%�U���lw��@'�c�������0���R�J��2$	8x�s�\d�S.��W@	f���{6��{�ƍ�0I�0rMFm�߶�����e��0I���j���y���eT�����=RP�#��J�9h����?$�G��GVCKVn���2VX���_*�xo;J`��/���U`K	u�i H��A4$L��r#1���1T�蛐��KʗB�@�k�ªn�E��ft���K�	R��t�=U��?���sJ�$4���Z%�dV��<�"�|8<�z "O`�5�|���-P��O��g�z.kG������C�G۷a�B�6�Wu_9`����p6���U)P�gi��40ӕ� ��:�CjA������qD�ࠄ(J>�\��m�Rj��@�p��8�� ��U����%���l�x�M��ccp�`PC���'Zm���X��MX��XC��Ce��&��P��Tb����Q��F�ظ2*�����BC�M�ĹU
��g2$R�N���������+�|X?�������w�c�Τ''�UJ�D�`l�N�~��E	��[6�E*1]9���TZ���C�y��{p�Jdb֩�\�>�|��7��AҘ��EYQ��z�$'9�e��b��d&H.}B��T���[DܕB*\�*���x��&�T�9��XFJQ��م	�H�d��8ǡ'�.���uʲ�*`�D��w�F �P�(4@�#��sqp� c����P�����Ҕ��Dޚv�9�	rY��v���a=�Kن���҈�����xg�H�E��4�L��\���qBbBnަ����qbEn��^�\��<j�
<V��x"d��Q	D�3�ŭ�Ҍ*I$hn@��0��=W�k�܈f�^^ 2������;�mݗT�	"8r:�ur<���d�$�`u[��H�ZI$CnU�NTx�����Ů`�	r��Qh�.�Ĳ#�Uq��bjY��)
]&}��4���hAdT%؊rX]!�5�����G=-b�24h��D�*�/dT@/��R q�iH� �}!�/���%�+q4���A ��Y�,d��HBj�e�L�
�WMH�;�2�+N���E$�������~��X��I]�t(,��:T�Q�fB�EP؆�A��L�1�K*z:ۊ��(D���X��D(�z�Յ$C\D?�}�\�6
�OJ%�C=lG��;v}u5��� �l�P��.C�N�3���JM�5T�U����&I������@��у��+��R���U膭Q��	=)"h�+��_ڪ��F���TU�y�q*��d=�8�J$�PS�t�g�9Mk9�U/�(�g�0��z7�!,��,_�h��Aڏa7�kS�E�P�$��Ȅ*I*h�P&��Q-H�$�����(��v�LxU�ְ��D�.Ub7r�')���4�Z�d���K@@�
�eh��Ɇ�|�pl�(�](e��	Z?E���f�/��H�L?�|oP�x؃��0`}��jQ���'��`g�Ќ�f�7S`b�J��r���3�l�2G�B:6R4'������
���<.WD}H�%J8-}N��A�1��)L{���=TX��^g��(���+G�F��F�uD�G�(`�!@I̹^e5�G��ij@�l�cZ�a�s�����CL	G���޼- �(e�ڢ�!%�7$�_B5���ʮ�	��;7�b�T�,Idf����yt6I8l�SaU��Ӿ%��F�pH�3���sIEC"����K�[�� ��Z�!�/�bRJ���-�Fx�"�u�+��SE�*�"T.�J Џ��N�-�+Q���"�-D�|�B�&�>qx��$�@�>1���h�}�R��#[�Q�A�Hzyz�i��)���Y&��33�k"y򋯔_����}�zD�;�"�����ꮩZ��.�,yKH�F��) �sPE�%CU	ly��ìb�H�UUTdj�o�R�.�M��ٽ��ƎI%1��bMoj��	��!k՞Y�m��4I8�Ԫ\�6)�JI\�ā&��v�R�cj[b�; �M�V�(�F,��<4*c���P�^�P�\a�d,RR�6|����̴�(�'��8����>n�P��!R���.~��w4F�(��3��G�yP�\L4I<��T����w.�0��2��e�������c4���B&�Z�ȓ! ��u��z�ٚ���ns�R{�T�b�yA�^�%��fkM
�L
���5U�-�4}w5������΅�Y���*OU�U
�F]^��^��x����SRUS�9~���1T<��GR��"�x'L��`Uܑ2K���n6��5��k
���X#0/Z�E �ĺ7PŇF�j�T��6�tAZ�
U�nRm�vm,- ֮���Hg֦Q�ﾢZ�%hT��Z�I�D�4�3`4W�"]i��|[�����+�{��� ���'���vڭ(��H�{�K�(A�h����@3�Z�~���K[+o�5�b�&��݌WCw��tO|�v� ����B�����d7�Dɲ�EC{k�,r���	�,.�LJSڏd��I*���۪|�j~9B@/��`����cD�`�ɪ����G�Ƙ�U
�C�J����}ޏ���wH���KY�vi��^����:�?K�;ޓ��H��+���������D���ĸ��*,ȌZ�`DC݇T�m$�DNR��#s�)'L�M����OG-A�M?��£��l+8�8Eblu.H�0)uhh���.\f�%�GM�f�]�./��(���\��#"��	�th��]`�������b~�>�?|>��¥	����
��s$y�_��A�4�o�o2�[�T�� X(@�؏Ⱦ�t��TK�4��P8��G��NgyxC$CoN�Pf��C4�:�%�H006��J( Jh�e.���#� �\�	7P�~����>���?k�+O� ��/P����Z_�q�p���.K�-��%�1)QN&���*`�
6�:|fM&���
��u.'��R@�V$	��<�4�X���8��I&��G#�F#p�.��\�4d=�+� �j�	L�G�jL��B�.�+��ֱɦ��3�DCB�d��#{��I+>�y0|�#���t]"�4 Y�2O�2TN�3 �J8���E ���U3�J|'�{D���g�2oPؤ&����r�Ƭ7�§&1�`�Fp/x(�p$Yh�/����L��W�1���w�Z⩕.�%�I�<���Ł02�$�lc�By��#U�1YW������Jh�����B^P�x����IU$/^�x�k���BOɋ���ըCr������'��E���D7t5S��ȭ�G�I��eaR��0t#ƪu�J�A8�@�4xeSB"h��F+Fढ��¤���$B��K�֖Jʄ]\#{�2"2#�M֐ڻomq�:��2�򍂒(V	���s�c���g�z��,�SMjH��C��O��_kD�C>΢��>���ߧ��9-W�.A���`H6�}p��y���<3Ɋ��!���� ��*���i7��Y��
I`��8��{,�,*-��<�����pJ�TI�Є.�yT�&zs�I8����eկ��՘C>L��5*R��+� ��A�����f����@�8�κ蓺@Z�\��`'���U���-1&��DvZ�D��֝�ݢڵ�SL�_�7eCX ��,UG3.����n�c��ʊ��� 
@P�(��  "�"�6�l�S�
�]���Nꐦ�B�A"(��&�Qp�'�Ks�y� 1!��k~)�zn���g�Ȣ�:��l�X*�~?�_��n'��{�����	�� ����{����������E1~��t�JG��_��1߱���a߿^q}O��/~���TO��������y�YQ�������@4֝t�Ns��q0]��E�p�"�&�MW�����r���ٓ������;\���r�gVM�������5x�%�o�3]|s�I鏮V�>�6`���;0�}u(��lG~DO��|��/c�g��ǣ���~����Y�<���y�w���U�3�;,]�o��������ܞ�������Ŭ���h�~�ğ����~/�&/�߃�a�����M�w�P��3�����V+
�<`Wy���_�~�34~��͑�*��7��������tS�����F�?� 8� @� A�@N=����"I`�`x�ВB�/���ʀ�!���C�oA|`�(	 �O�1v��(��e��c��|r���8��M���.����h\X�����oUL��x�ӌ��Id0Ybk�K���"PP6;l�`xV
)*Ga��͇��;?��dDʩ�h"-R�=.�类.�����!L�����P��~�%7��r��O��Ny���>�ۼ��~��d;��箟����� &�`��y��9σ���_�7��]��G;���!���'��j1�C������~����b%x9Q�����O��WӖ��E�)�ǟ�|MNf��m>F���uS�h�>�[m�>�ޑ{h�p,�h�^�P�F�������E����OC�^�^�	�� �qV�x?A�|gE����t~{�ߌ����9���N?���~��������m����"(QH2���ߪ���%W	���@a��:f�����ۏ|m?���?��o���o��|qϧ��！�ג�q�H���g�ɍT����=��<����R@ $A"�"ڋ�Ru!�C�Ī\�p������C�֞����3���?[pp�H����w�J�1{�6v5h��m,���'Q��7��P�����d���?��q?��QLb��*A��� ����W�Nwl������,�A(���^m��pd0��?��~��'1���~ި�76�BB1GZ.������yɰ'K���`=����>M;77��{e���x��mS��},S���k&����������-h�?���]���p`Xa��C�|�3k��g@2� e��wz�!pqܗ]��7n���'f�`W~�����B"��3���n�+���>��u�!/ϩ������y������'�}k����?cn.�ψ� ���G�h��}�x�wr��JGR5�_ζq��q�w��4��@�zyi&�wp�m��3O�W����PzO9��;�, ��xR7񼽨��J�	������\���n���8���E�}[$�$���8NO��8�vB���'�1?����d䤛�yP��#�{��+�@�i��N<f��/澕�  HH�H�$�� ~�8?�}rb���d$I �$A��� э�%2h�4k$�L�+(�`�O���>�ȱ��<H��v���'����3��X����5!�����"y�8�=�:Kq>f#��y>H@��d��[����ӂ�u6�~���AE���}�j�����}�g?"!������#���n�F(�m��[x�Ů���]7+��;�9��E	F��rwrr�:]9�wr�r�n���w:�wF�r6�F6�l�m6�Z-�`Ɋ
�c1@a�If&H�,A&��3j�4���5��/q��UD��5Qە!Y7Y�ɦ��U!&�ƭA 0p&ۅM`�ɤ	��%Xk�2�$Di�kU����ET��I�d���Ə� XR�
S�#J�!�K�͔a���DF��!qF.MP���W�����*���i�.�V
Fm�HJFݳpDɦr��OfI�����������#$a����ɹ�>���,�(�r`LD��DJMg��5Ģ:s[ү6����k^�z��$�IΑ�2��r�����s�S0ƅM�[���}����*���jy��2�|���u�s� �̙˳����uۜ��DW�r]�!s�wt\%���U��ov��;�Qgt���WwW+�+�wv�V�>ch�0A�U01���d ���K�h�g1����pweW��۝�ݹ!F����.�8�g	� �U0X�2Ep��.�;b��.8��R*( i�����Ҟ?��)��r?S T�~I>�C~�%� a�TZ��@�,a�!�\LSbF%�|{x��E�4�ܬh�
A�H%[m�"�P7yn{��r�"���Bs���B!D��Z�E��1��#nZ0&PbVJE"F�`ؒ�@%l%0�,h�"��T�H�� ���R�b93&L�ɿ�3���-FA$"Hķ��l���6�YF�20 Y*�F#  Z���s�QQA*쐩$����T U��z�*��H7�Qk���!#U	HD�Lr"bdV0GI
��U�s�����e�x*����.�066����_�x�ь�@>�}L�M2�?.zέ2�`F�%!>�}�w�����ݳ����I*<��1��o2K\\�$d�ں�RJ>Q"D�l d�}7�L_�����4y��ֶ��M)�O��3�qϯ5ȓ�6n?̘�h��#����c	;q�l�W>�)4��q��'��~���3�3%�n���_xq�?���UR�F�1��$jLȆ<X�m�鬗��I��%�|���=�|��䑡<$�Y�e�'�ӳ�d�>���#!�3��Ł@"*�Z��P�pD.!༹�����!s�x؄�(4G�.��"��B�U4C2tG>�W	 �c�M��ł�F�l�͠- ��A
��
6�s)�3bau-��8�i~�x�M�g��m�M0�e�& e&���8�
���y��A d/��c�@����o�>�iH}��!���xP����<<���X�n"(O��>�� �(�,�C�6��`�
�>%E��e�j���b�g$
�]�_G$�Q���Id�c|u�>���L���c�����c����գ�Y�y&����0�$�9P�� ���㧹�l>�,}x	�߆�o�kc.g\�W�.m������d\�]��s�7��d�����v&9����eY�XB�}��>W%�W2��|���Y>o���	��,�Λl|�����&�i�K	4�τ��!�@��@��PQ\ b	I�!�|˒����$�dǈ�5������8̺��6��,d�(�"ݎ&2X�ϕ�2�ɄB�He*Js�\�.'�a@2O� E
)��ϴd�J6�hx@02�RR}�g���"S~FQv�ݸl`j��J�7t��j�-�|S�]�}������3Y�#b(ѣcl�s��ߴ��d�>��f�������T�  0Wi�Z�8�3a���w�x���VwR��iM4�	kDL������XG��I4+	VXi9uĺץ_�7���"�]���
��`�Qf$�@A��-�od���s����t��n�	����	n8B}�3e>���{�s.;&ݗ#�f-�d�>M����.�D$�c��1��Y7bM`i n��@�w���"@��IgΙr�%��2kj`$���On�~̙�$��L�h�k�Q���H������}H���&�c�UB�H�U%*��jE�f\E��d��~���d̦C����� �(��*,	���������}���-�}�ܤ���h�7-A�ț�i����ɊHI!	���LY��(F5|����z�(�H�BF17ٛ��5�Al�\��r��nm�������AE`��PP�$`� ��THl$!,�������1,��`Q�>�C)�"]�I$�#��" P�E3��^���0GI�BJ�Z�z�r��]�sTcUq���S��z|�����uj��H����r��BI!�x	�NB��:Jc�!��F�#L�61�BQ��!h�����]ۜ;�� Q���Hl��o1��3����z�h��!x?
w��	����*H,��4y*�E�RD�3���h�DLL!�
��='���\~���7�3a�-j�ZZ6���"U�a*��Qk2H�30&`�lc��jX:������v�s��n�� -2e�I��D�qdTQDL�p@�g���`cS�~����	J���j�'�(yx��G��a���U[&q	�R�*D��8߉I�A8?m��K�2�I$$	�P"E@��:��!@�)�1I�D�黗*Y�8����^d��m��f�,�@�)k7��1� H&�m�̟����~����Dc�?��+���;ܞ��4��ݤL�W�t�B�r&��j,�s��>Z�#����T�K��(������[wІbwv�m�6�@Q'�\T�Zf(C��M�Y�'�ޟ�G�X��+Ͻ.!���!m	R���Hi2��	��#���� Y��f��Y�[�Ǘ�\	�xI�O܏�f��Y�k��7��qL�/�Ȥ,��Pj
�ɹ	S�R�[d���1����Lkǥ�N<�d$���0ə�M�߱���L!�i?� ]��@HR\�8A��8�� 
��U�5�U�QU2 mQ,��_!��x�٪b�2�! za+��d.�� 	!��i������re7�����n���M�}_㯇������_O���q~�~���"�:S�:�Q(wc����~�x����t]׊�7l\>��ܽ'��������9��$p�����_���W���)�x��A$/��}'�?�w��(���/����K�t�&�踱���yQ_YĿ���G�/���إ�;�Ѱ� @ A� 
v�A�̛׳���&q��PE���^S���T�$@���P�A����OjAq'�J\ ��UG%�xk���AGjtH�}E��󛵕2'��	�]8j���j@1��P�d@�V)@�N��F�r�s����� F�Q�N$i�f4i?�m�J�ʅ;��
#�,��Yq濵�I$4r�J���Q@~=��6�!�(�H ������
�.��x���2�B!|8|h]@	�X�úJ9�K��[!y��
�DR{ďG��PpR
��x@���# QP�ŉ�8l�/m�.��������������~��^{����f������_��������������6/����e���ޏ�o�<�����?������?�o����G����-��I��������x�o�b_����dG.O��7ᥱ�dB �����P%c�e�{@�u�e�]���Wn6�HUJ;����DI��� b��kJ&8D@6�ݩ_�t���ɱ]d������Ó����A��������	��_���~��?�z�������l*s�Y��.?�F:��t���2�+2�o��f����gQ6�~;o�%{�q�;�h�aMg�Gp���F�d)����뮍�M�#�׮Ъ���n�>a��y�Ma=������D̻V�ۆ�R��p���q!>��D{����TB���Ĉro%\MayB2&�^���"# �I��"���a�4��/\Pu*O������ }�	h1b� =��ϫ>�k��b����d�`b#d��*�K( T��P�w�I'Ʌ2\�\�g���7.�y�����]���ˁJFA���C�ׯu��I�KJ�*��*��!��$�d��}`���+,g���ʻ@���(���$թ�L�3��C=���U�(���`1|�A/0E��Ƙ�B�cċ��!�	�ZI#!�"���/@F� �"#z� `�Dn�p�-ʭ�`H��/-��8b��}�����C>���1J*�8%�38�O��v؊uhU�4ꔻ�R����s �J��nX�&`7nK	��ӈ� �4 P�P��qP
�s�q� F�L�v�+P&���!~����8V���=��k�x�Z�*Bִ���f2S&�)������.�N��	�-@AQ�u���@�p�@yr.Ǿ���"�K�qW�R*+�m;���D�G;�\�����с�,	�~X�h�F;�5Ԋ�ٰ�`^��EŲ� �2,�$�� ��
h�Z �&�F�Ѫ"`�}]�CF�51Hn�_�~A�D�o�](T(	�$4�D�BBQE&C!�R]ܖ1��/����cQ���07b&��v�3� Z��N�b�� �"9lw�[x���9�k��(����pM�H�hX[�w��
~�h�4[�q��X[����嵛%��+�(��K � ��b-�@�Bw��)4����7+�Eo�F��6H\nd F�0�79�U��,uҢoUA  ͍�u\�&"Hg8*(%�`
*v�A�c�)��ب�`�UA�� 7�_n���H iL��7�C!��&D��$(Tb&4�7�[�Ƨ�UsU�Q�Nqt~�`w�8r��n�Dбjе��*�4]��)� �����*g�#D1�.p�j�"��
�!�����۔�2��� Cb���� lbǼ�c>%E*-EdF�!.CJ)"�BF� �Do]�@k�b�7B�B�Ԑ��s0�,��$ ��Kk��-

GqU�pmܰ�33?�֥��0�DA@�@�� `�0X9��������$(�R��{�ל��p.y�~m��j�-�lc.��"W5�mΉ�s����U�+����]s�wnV.�61�r��]�6Mj6$خgu7qrd�]��I#!�dD�dd`B )�P�B�̹�8Ӥ		 �]+r���t����15H�@�*��L�@�i�5Pd�$HA�`_A���@ъ��R�Utʠ]�WsSN�ȯ�)�@�N�p�QLŽ`d�[d/@(&�#�y̼3�(�� �ρ�uF�"s ���>��(g�]3		$�]Uɂ�?��%�M�AUY�֑՛��a/1��3y��>w>��P��f%,E����Bpn�!�D��MLU1o��6�ɭ�� �XjU����oԱH�C��FPn 0!��;U�Į��,�udV�@���E�tU���&0?­�qU|�B�$%5J�ʲI%��`�qp&@ 7��n=�\�s�GDl���/`(�����҈,bB�b�#�R�)b�0F�A3�ߢ�2����`*�� ������!`RGEL� Ɔ��g��x�Ol6��H�F���!$$�J�@���E� ?qST�<p�{�Q7�{dX���Rj�3�B;����l�\���. $�&0Qtˑ���TaW�~���s�n#�P� 
�,� A�	 �UF�A �[��O��k͌!$ Dd	 $dIdVA"$D�TWǸ�qj%�K�ڎ���{�"��1 ��C⯹�?�>�M!��F_5��w޿���!wF"4]���@9���r���i�3Zf� -׷���#�[@��*+���m  	�"�����*� F��pnm��[!�F,\��(�W���X�@�n`]�����9�$V ED(P�*�o��]%���oҩ�i4�3U�	�%ڰJ.6)�
5Ɍ!�d�l�6�8��?,۰5l�[J�l�����TWvtF�U�F�ͦZг�!�5����1���J]�L�οG�a� d�СD��l�\�A���x�AsTK.�x:0��ЖC8����Uߑt��^��ʚ@�!!t��A�D�P�P��
.�jj{�v狱��,���zZw��l!�W�Qn��]`��;5���Z��F%�@�XtI�2;r�����9�?~3�����Yu��$1
(~_�P|�4 B�q)�6��kg��Wq�y����A���i�!o�z����_��3��Xlm�
���/������l
����Bo�<E�_��~���O����1��A���xDH��O��@D��-�(�A�R�IBZ��4k�������x�����6U�@&b.Y�Pt��23î�i68�E s6���a,,ɑ���2Mq��~�	�S���h�Pa>�� ����yB�	�@"-@����@̤�##9O=�5"ᄥU�_�`�Ȓx��/�g�3��� �!����b6:�D{�QI"�>)��ӭ׀��o���	A@�E�@��� �I:Ǿ���@B��yI�$����r��UR�� .^7�Q9D\0��B���O��n" � *�(�?������u��n&��I�Љ�pW6`�҉ڔ'H\��oڽ�$]�5��xc`ԽB���g)[ (9�M<�u�ڸ�S��{�:G�0�.8lv4+z�B$U$A���NϿ�6�,�<2�������6�Nq��P�ۂX��H X�` '�?e%��B�$qy_�p�xHX�@b��>����2JV�j��� �(���4yV.�6G����p}�����ⱔM)Ŗ7��o��( �C�(���I�AI_w�m�;�:�V%����$�{��"���nl'��fCӰ������q���ͧ�����O�o��A~� �BH0����,�!ɽ�p��Y���E�@N�dR�H��UN'�Cʱ��񯛽�Q��"����ı�O�X���@��$��6�� ƌTaY Q�@�y���p��,&��#��(���F������P� ��  鉻����Ha���|��ޯ�07��\�q�@�i��~��5ǈB��O4utEY�|��O��J�� :3�B���9�xu:
��h������hdO��
������&�%�V@@$PRxҗ���RwI�R�6��g���5�_���]�7�Ӗ7��Ǜ���,�0�Bg%
g�/.W�q�-���?�aypR��lm	%�zhv%�?c��d$x[
z�>櫔�z�]�<ί._[�q���@��;-G���s~c��{�`
>3;�~?��;�����5�9|�����wO�{��z��@�|V��k��_5�����C@<��;i]T�7>�(?i =R{"��g��B�H�@� � (2?�pa$#�V�q'�O!����^?_�ږ^��!+ a(yb � *�<���ٹ�Ğ���@��O�x?�-��.���������� "��(�oA��=�DB����	9T�_����L�¼�C��(JV��ɾXN�"���ߡ�dP! T'��;�siʾ����C�1s�PܲI��t��!!�x�. ������ !ս�^��[3�yl��g�l��������W�P��C��������<���,�G��&�A�Lv���s#F�K��?�2�:;D�����C#6����t��|�F�"����2�	_����*4��4I"2���<Xs���>�k����>ǣBJ�v�.�)N�`����Pq?���y��}/�	CG#��X�b�zd�.��q�JA�Te^�Q	P,fa����hj�q�-K��pk x�)B�%�C��j@Uō,q�Qu����*�i�a����ҍT��-����_l�*@�a�0NW�D���"�n�w�u�}�������k�Bw�T.���os!Rq�a�C����S��'�������>��{?��d���l3�/Ql�x߰'��0�}G� p~H�cK�����`#�����,!\�G���|2֭\Z����=߾�>�����+�v&_��g�;�;��\_1�?���5�s���Ù�f��t|��������_pS*��"��s~G����;�Vcߩ���|S�L�Β�ߌe�c�IU�3��qc|T,��G�S���MR�}��4d!`�3�F;�/�J��/��78��_��Ҍ��� v��(+�z����������\쏡�A��IS��s�����@� ��U�ѳR��:���	��K�!C�]0�����`�8���/�~��?����o��/��+���'�;�1)�d�����Kv�d���LOjG�_��,(�����c�2��,v�i�3�ߙ��ڭ~\<	ɐ�����jN�J*�A~�=��?����/�>ֻ��w�(����! ��a�a�]AG:��J?O�2Ұ�����	�c3���Y(�O�F2a�R&��*u�")kw������@��~z��X\���6B�q/*��#�6e$�fX��k�(�) �T̽����/� �\�W_���")�Jѷ�:�V��g���R=}���w1��ӽ�N�k�1a�4�{�9V}av�pr@��z�������3�uE�Z�l�$c�]������}�~y�=s�@��"BI.֛�����ƒ���;�}������4f{�w��'�8��o��@2u�2K� ���}��>_�����]���)*�!V��� ?�LfL���N,)$��7�	%Å\�m(N|�rC(C<j�Gk�
e�f��u{\�V�Q��)�;�T�9lG��$@��aJ�� a�NO�ӳ|Ԓ_�bg7�Ԑ�f��w��l�垛����1b'�BI`������8�Cˆ0����BC����(�   �	ߔ�풀
,\(7�2�>��2B H���a$Љ�T���I,�y8��l|�b�#4�b�i�}׾�W��i�m	��OP�{�&+�y����[w��9��p]�}�;��*������7��[����j���������������O�G���_�?흨{_�+���H�N'�$����;�׊�����{���_�q��1��K���$"^ؤ�aU�/��_�6� ��!/�g���<q�Q����ч�������_O�~yO�mn�A��e�����`x�/�s�?P\ t��pw�_��?�#s��ؐ=#��8aۡ��	˄�����!`̼��!$�,'��		G�iC�D>��]$$>q�(��a F��ڔҐ��xwT�y'�X�n�	f�'~���� � �'����!g�Ą&�.>��̞����џN�f��B�1QXDBD �X|� A.d��jA˦I%^��^�M����R�����0A��V
��`�"�(2
���tW T" �U��ï���R}8;n���@�{�a��.!b�"�U��R*�HH����!�wy��EJ"0B !�MDo H��Al�H�~c���.C]��Yw6�I$�,!T�R��`� �1R(R((R(*��y����#E� �(���l�6�8 b ���"�'�J_Z��$����D���V�ڒL� ���@
`� A"�P"��� AX#H)b$�7�Z,�y��7��E�T�pTB�(H ����UT�	@pb�	$��Ͽ���G�ĉ�z��$#c(���@`��bI�����o����tc�S����Λ}&�[���q�X������w=�{������W�����ך5��$���םQ��X��HbRDP�I!����4��{�ɟ���J]»dR��1#d���������ݬ�h����`ȳc�D�P�v(#[��в<]��QFu���\��S�0�3���dL��;vbi��۞� ��'�OZۈ�Cnu�U�a%�K����J��!���D�� �
�b����� (�V F�P�  ~���\4�hJ�V���􏜑hY�Nw��������{Aj-�mYF�8+X�v��
�5���LE�s~�B�S�[��}{R�h$�T��X�#I���Eq
9�I�)P�Zs��U��"�����j���gL�}���_�e(�%<^1�n�����ͥ9Yk
�&�V�cg�5����XZ��IFW�"ƍQ�o��8U�R�@�?�)Ă���ADh4_�l��%ח�A^��/�CkN6Ih�e�_�.��6{�ǈ�����Q{h�J.v���1HZ9ښ��i7��+*��b�JOV��D�T���hXSZ[g�P���4���|W(�P�Z�)��&�a�4�D%\�B�h�-�k�I1:�H�Z�m-��/�R��&�km�����P��ii��ڶ7�y;_cg���d��t��.�թ�g�TI�Ka���!4t�!�]����g�FS��E���E~ᣣ�Pi��'�Ʉ�m|�6�\�L���bD�h"��������t�nv��?��5������Nt�;�j�աH�#%��]��ۉ�|�~�R�<C�r�k[,!�[o��U�s֝�l�b5�i9.y��2��k� ��/�t\���!�s�G���f:ΜG�鄌��i���wI��ԋ� ֶ��J�����W�g��^�M��Z��l�'l�}�u��/�)��u�;�4IF��jm��2c)Oq���6�e�1M�ƻc��E�jN�հ_�vޯ����]=i����f[Y2mw걣��Ҹ��+���
uȕ�7�������5�j����cQ��ӛ�Vw�+�ם$o���2�2l�PI:1�8����~p�ƹHu�i �׭6\軤���5�$��� $Q� �j/�m����O�q��~�^���GӍ)�p������R�kos��6�c�f���Z�=Dw�k�H�ݴ�6�c�|S�������s_^��~!��d暴�%�����u�@[bٯ]�ѩ���t�f�;sW�^�A�6�qn���Ï+/7G���n�͢�q�Q���],��+M/�2�^���q朊mO5�&�<­'��En�C�;_����4�1�=��Ξ8�v�t�v�7��k�j�;uϙם�i�Z�����~�C�׍����9ϝ<�u�8���8��%��o�|Q���Iw��9�=��{���ΖK�������۴/���|�����8�<��}��<��;�3�{ƙZR���^�?/��(��F�v�q���e�������.�g�Ϩӈ|�qyiZx�@�]7�����9��/���M`��   �\��?��j��Yk҄I�M��@�D"	3!b��S1�T,��H)H)�)b,E��@���|x�s�o>{��__^ϕ����q�&<�?}���m��O�m_�~:�p�7����sGI��N-�R��ΗG�!��/��af�l+������|wl���v�X������޽ȯ�#Eۻ?��c��hq�5���2��wϷ���֘���|k���������~a�=�>�}��4Jv<b��>��m��Pv���onޞد�����'�~���J$0}7^t�T=p7���7�Á�,����}:�<S��~��7�f���Z���g���1�[�o�'�#�
7�O��c�ÿ���{x�}����Q����f�k>1�����ɷ������t��<����\{��5��g��v��/�kg����O4�}��J4�ox௿\k��3�/~��O��v���ڑ��/�*޳Gq�ޫ���n���~�^�����o~�w�K�T�Z����������hg�[����~��ϯ����~��v���Ǵ��4nWJ���{{�����Dr� ���88 o�����/�o�eͽ<�o����|S�c���9¹r��6�nF��6�Ϧ��$k�$��M	��������TǤĻ�o�?1���A�����[�n�Qn����G��|�y�O�>>sַ�P�lV��Hb7�^���x��#UX�m�N yȐ�1�iq�C���z<��ʄ�5v�������{m�O^�l_۩o�>���
��qN���6��ô��|��:{J-����������==����=��Z�{�宿_�����߯o9��ޝ[�oOc�u��������]4YX�b|�P�ô�E�0z����	6�@��4�!G\�S��sV\��M'GIq�b&�pa �ap!��h8Je�׉8�4�a�!�1]UvZ5>2��Μ��Q���𞄷K1�\�؁1!x�Cv%$��x�I�ޚ˿��op�o����<M��#����F?=��5��0[���c�#C���' bͺhA�m�B��b��F�4J���������6i�~co�x��%�w^w�����������u��{c���
{�oqW�د��s��`?��p�Pu�����U���Ӓ|��'���	�Dk�k�����5YV91���Uy�9�MW��V��&�BluǛV]R�d���k�yU�\�ɀbPs�::I� ��$��LD�\���^A�I=b,8r¤���Qq
�4��h�e�h��RC���m`A�<q%�D8�d�����4Q&�1�FB�JC0d$9�H�B*a�r.�!L�z��qF�΋�(�eNK� B�-G�5׈0'`W\@�a#t2`wDH��]�c��	�7Ux�<�^23I�bh��.
�8��Q���e	$��KL��(�@C�:E��9�(�l���|r�����&J�٭�B��,̑9�Ĉp.�8H��?/��(Z.�3��l��!G0i�a!��^<YcP �X� ��\DN�N4�Ȭ��Bp�F2�7$���=$� �LA�5���vh�ӊ+��K Q�.�0��Ӱ��L��
�(�T�
�.�F!iC�S�M�Nc�(��XY�%��r#�zd]ɥQXH$CH#�G��a�L��$t8I�Xl�R(T�`��xr�lG"$��20��*r���)!���.jΚ���̎무pN��!.C�"�MDG�	d�]��7]�Q���Eug0�6X��nwBv) ��Il����������2���3�%D���Ph�0�02"�DХ��;o�N�]����<Bf�H�y�<,oP@�Ǐ]����� ޲�HQ7N�44SD��x�X�)�*Ǜm�7GA_!�Ky�ݠ���Rv)j�5={��A0\�%!T	�y��.Ag���"g:����*�B)�,$�I�ؗ�d�rwq�4I�D9aĹ�^i����8�')�_�^�b�>Y�*�Q����UY�8k�6O��sYF���R�u @�J���;,
��P�U"2�`�ԣL����F���p�
u���\
�Ҥ��S�PJ+I>��ZT��#iW%��*F{,��V�)H��4����d��~hܜ-!� ��c�>�e)�T�{R���Q)�c��Tt\�C�"���MK3�À4fP���	�t�'hF"������"���C����OM,UEA�t�\@�2V&�M��,x�)a���5RB@�H�3U47�hQ%���b>��FP��lSʱ��QA+���X��넚�ΐ+��zqA[e�3!��9*B('�;%9�DS��i�y�@y ������X`��f�U�f���Rt3�-1A�"�@��VQ;�\�T���	N����1�`$i�#2#���$pQX)���g
���z�5�TL���l �!��Uy�A�)e4�C&$j"��J���Q��:E��%&^!�y��>f)YV�@kД���JN\�&��JÇ�����㵰��QDR�bC��V��
&�ل|��xﱌɛ�Y��2��-���K������}��U�E��0B(F(R1XD AH�@  @��^����,�$6 P�OP�D������OB������P�*�`b�;l @�9��*��b��lk��q��2<�ٯi�C�W��
e�iB,�'y��${�t,Q�Q�I�h��Q�T�M��/bDK�Yd��5��#�3�Td/��%c�@H@kA%��䘒6�q��� �)/"�@Nv��5&���d�C��/;)�\�/F�%�@�Ҋ�K��jȆ�GM�3D$�2@rEx`J.JM��(�[1�>�^
G�|p�X�<��1gZx�]up@X ژ�m���&h �YAB�f�d��ukk�"�B���`1$9.�7
����%
&z���wQI5�z!���>��JKE:�^�Q�p��B/�d�ҎL��F���b&˨1A"5���/�ߦ�8#c~��2���Zڪ��T2��n��U�d�g\��PU�+E�|uk�8*�3ͥҗ$�E<i�>�����J(��2͔�(^:M@��i�h�)T�=(P���n�H`�n9��(E��!hR8�V��4�>�C����L5�KȉU5��h�
���;V�[��w�9HKJ��26@��&���M�	� ������|�Z��`bИW�@����	Eb�!�A �@s�1��A�OxQ�w5d3�
�o&�@���:`ԜRK��"����%PQN����#<,:�K���Z)��v%�M����W��G6gڑVxj�Lp�n�hprIu����0�<h2�ԍ-�0j}FĴ����Ke�+��JiBL��8���[ ����2II����h�S1��0��􃷼����g�1/O�Y�|)���.��]tO��������CpT�EYB��km��mۮ�����Bc�����0Ox�A���ɉ�5WF��g#F}��<�˘AC\���;��Ұ�S�0}L*�n�g�y4`��X$��+əKQ�a  �I�Q��YjP�PĐ�U>+ZM����(��eU5���faL0Y�] ���
&_�����[D\:§YSDP�Ȅ�B[	�J�q嶁�J��sg�D�E��x��(&��UV��EjN�i�'*U�����/�̣��)A;n2r
U��\(�V��%�AY�=z`A�7b�������lLU��+�]��������T��KKJ�ew����	$E����?9ҙ��4x(@�:Y��Z h���y��,HN�<18�q��,1a1Ж�tJ�j����=�YY5]И��/Qj�a,j�tQȴXya�JB�_�&C5r���8�lA%k X�u���f67qA����4���2�F�2���X��b�X�q	�t,�;��0����'@n����(�ވ� �&h���1���.`���5����oB�5�ؖU�j�&ա�;�zG��,�+REBi����h��n�a�D�R�D���!�
�Lf3y�Ix�=�ˆ(��9�\(�*��n�<ӘcN�
������2�`�	FW�`U�Q��Q�sGl 1�ţrG ��0D�A"|1V&*�-��� �8'�.ˍjc�t3�1��AHa0�B	4J��@��E�K� T�����ו�<���ZwDt�:\��]ɲ4�D��L�esº722�T�4DV��3H�,&s�eTqטŒ�H@��V��:�.3*�P1i	�+�1�<ݖ���D�0D�0�����K ��4(ja��6jrp/�[�8u�Yc����l=���q� T
 ��"5z�����������W�� P�,�^~�^�kmd�ߔ��o��p�/�q=q�jRg��2��K3���1}�Tr�e��Z�Qť�ψ��|W�(���U�������M�Ȭ3���5�Լ�j����+<��4���Л� '���p�s!2���Pس ��^U~�YR���&�܉R������ �����2c�ɱ��$�e��!�%����Q�䥈mݢ�ա`��'.K��Ӯ^;��)x��a���=�:��ܴʨ��&�s����Ƙi�,��0�c����vr�ҒV#6w��N���g�������^�XZ��^�O"L.ȴ�>�˲�l:�c�T��]x5-,���-X}{Y0�*S����tr>�H>�l�F�Xx˙!�K��9�:%њ񊭢ɥ�Ӗ$��TYt��)��Tc!Rc�\+Ń!)jbg�����װ)m�'�[R��V�<����!XM�R�t� ���;Z�	O�A����T����Y��m̱������)Z�"��{b܇*e��r���b�e`a���b�DH	Pv�cp!�:%m�����8��6F����Ay�ƊP,�5�C�2�1ۏ8��2�P���(@Hd�0�ڝ�8;α���O�T�EV�AM����j|v��-D%Y�Dhr��̾4��[�3����̾,���������c=� ��J��c0��z��v��6��i��<rrl�Z�ۈ�1�.'�=�9(tGY;T�pZ��4����,E� �j\Z�[(�j�h���лՋ�>p��1�y�b���$ku�bU�/�)Tu�&�4���g�����=z�:�N�B�$�L�@-�.Jv`����V�e����C,L���,�(:(�ظ׈���B��FYO�!E�&R�l�q	�4�����1�FlJL%��A��}������H�/�/C�ngّ��� J��T)E�����J�@I
@� {8 Z"\��TUD�A@�bX�*Jh�6ͥi���ջ[sFŰ�V*��Ŵj5���j���Z�lQkT[|UsZ5��Ur�]#D��D�R�o-��5nV���ڷ6�Uskk���ڢۛ[�QV�<���Q��[sm���\�-��Z汯���ت-Qlj4Dlm����W�-�lI�&�Ch�RZ4$�j�E\����+��;���nI���.H��{�& �ˏ92b(\Ӯt�+���nF�\וp��ll�%�m��lͮ\�ͣQh��b�r���j��65-ccE�0m1���ڃ%�61d�AY$�JŴU�1��CEEd�X6��[ص���X�EL�cm��r�b������*�k�Qc[��KRj4Z��Rh�dY!@�|����p�������ɦ�������=����i��{C����?��o�|�>��o�?��z�������oto�������_})�~�o��ϭ�?�~�����������=gc�?��z�����o�|��x�K����__��#}��<~��;{���������H�Q�CP"Ehh���h�����$���1HL�2��Dkb�%�f��fb�Q�5���E�QTVѴ��5�mjJ�i���Ed���b�1��ld�-E���5UH(�2!"�����HF�Xbk�HXѬ�-km`�E�$��E�+lXJ��lF�h*����l�UF*�AUQ�j�lZI �I@		$A$$�UII�[AZKD[F�E�� !"�$��*� !j*�kZ�6��������KQmd�#DTV5��l�ŴF��% RI�Ѩ��(����$ذ�26�EhՊ�H�H�H��) "�ѭ�m���kQ� "�ȈH""�"H�"+ � �ȨȪ2"2"ȊȒ
�"��
�������+"��  H2(���"�$�"�"# Ȫ�
���(H�""
ȣ"������ �mQ����V5j4�  # #"�H+"ȩh�mZ6Ѣ���Y$AdA	�QVEQ�P�AI�	d�EdU�BD@A$BEYd$$�dT$I	 �� ���<+� aϢ\\\� ������=w������������i�������܍�����_�����������7�?���������?�b�����������w�_������������Om�n�^|��m�z��������=�'�s9��x������۸�������?��_�������q���~��_��o�S�;�>���}�@�[���>ӿ�~��U�w���?�����&�
$ ʞS��	an��!5�L%C,��6)6S)�!��a��%Fe%&Hd��&b�M$�)�1
ɰH�ɦ&���JHd�����b�)�@��P̦ �l�Ќ ��BB�`�HbdQ$����B��%1�
I	Dɦ��4�&&1!4�,�,I��)�H$J�C �H�4�"FQ$ą)��Q"Pؙ0����@�#%3��h(Q4LJ�P�d2�K(���$JE�$̒3I4	����H�ِi�"(�&X�%262PQ��E0"�E��i��M&�10d��Q4J
0� �&Q�(��A��@P$�c"�I�i2�H�� �Ba&JL��DMHc#)JE��D�D�HIJC2a������!a��@!"HE�͐3K4$ĠJ&4D�l�ɐ�i�R�Ȁ�F[���P&$@d��AL) M$�R&&,ę)&�I�L! ��!��S2bc!!�2�L�J �e"��$���R�%�?w5��]��|_��r~�z�^{�����|�/��<���\������=7U�pY|�w�i����?��O��>g����c�����^��{�� ����85�dQ:ߋ��n���ݷ��>O���/��.ӽn��w�����<E�p���������J�������/�������}��/��k��g����?�{�q�?�o�ߵ����_VG��i�}��T�]���d�;�ؿ�v��^C������?u��E�鹬��7;�ϵ���$T����p�V�����7Ɨ�ɕ�s뜿�0�q������U�/����夕d_�"<٩��G��b�過�9(%�D�)3��B�p""; ���jDڨ�mG�{lOp*�"�l�.F5}�|q���"����X6B-��0M�����f����*W����"h��ϼ�Q�v�)MIg��͋�,S�^m�]rU=����v��l7�$s3xF�b�H�0`~�ce	\яB�$o2�n5��Qϑ�X��}���	h����ϞI ��Z���u���%��	lV�N��Tm��]�A[�`�IRL"�J��
�Uְ��>�m�#�8L�-B��D�GCd�S�A��9F�=��=���R�!�>���	�� ]�	�>;ő͕}�b����h���R9p�p^�r�xa��(c����B7Q�h+?�1��4=#�Nds-�kj�BG94�k���NbWT�;n<6���K�9e�8�p��)���4��2�UC
�b>�bP�!�Ub���7�x(l�(ӧ���su�U���v���sB �9�EH4�2���%�\�I��uh5�fpˣ���^m������s���,�T�M:����E{�*I��M! X��ˌ؂�r�,��3*�k��fk=��k-����KG>�\%��.낇Im�h�H�5rtt<ك��c�%��х��~�d��<��<��a{:
�K$��0��B�E*���e�a�9iEV{�G��a=�$���;K,��B�.�sMCk���QWm�n9pa� ��2����k�0O[��[�Z�|L�G�f�����`*�P�yEZL8y�`K��ᅻ|w��e��z��1	9dpf��9��6�_ �f��ؤ��й��[��5I���-Il �㙓oc�|�p:���@=�+U�b5�Z�foaF�D�u��<g`���m�L�*ENc�f�+Ĥ��~.ƢI5��eDD~J�څπ�*�g�+ޯAv9+�l�'M�g��k1a�C.�M��3M�����������T7�9�	� H;��?lK�|Q�ᯢBE�P�=TV�K��tZث$A�-��]r7��� ���.���K�6��!"�
�Zt$O�C,�a�Ԗ��%U(�_�DB�B�� d�B⾔�Q@�!��P�-Pe�m�����2m�g�����)0>|,T�D2E
#Q$�a�qZ��&0ǊŮ�2�v��#�!h�E�c�%��vL.$�7F@L!�ZtV�
]������-LQp�tLQ�An�ȃh� ��7�$/��)i�JɟY�f�4���>��)2SHE2K��r���
�b�`Z#h�qAr�*e@Y���ET�C$@=TT��1@�o���ĺ*�� $@L�A1F�/�Z�G2b7��f�#�0�gAK�����*���27�\��t�
_1�P��3!�8�a}(a	qE���"���X8]A�G&H7Ep�FةYK��D[�AQ-���*�/���T��*h�*��7D	1��q�rA��m��@mqArD�m�CQ� f����dI>��x�$�����T�-4sQWObAm���˗n����8�mջ�f�_�����)���Kj�(�������������������������������������. <�X��F�n���73��o��/j�4�Ҩ$��@09�8x��J�f��P� _��     �    �           �    ��  @               � �Ԡ  q�    �(   � 
����             #H@< �6�w����f @   ` @X  �� ��QJ)#(sמ�z ( )J)@QZ�B�
 �     �  O� ���    
  ���@   	� Y��     :$�.�  �    �%UoO   �    � ^���     � �                                                 <�  >     > a�    `>��8t(  @ �    U  D"PUPUD�QT HR��!B�  @     ( ��""���J��EJ�I@��T�=�|#�dK�� �%@���� ����� �@}��tMk )RJ �҆�>  a��/��$���5 
P�(8	6= �� a� �         >@  z��޸
@�� �0 l��u�  �  (  �� 7L   0       �  �)��:>C���      L 
�	������� L!2 �I�OɦTxaSCQ�d�yy	��4�S�S�y�jz���  ���h�!������� 6S��L�P42��y h  ����h��4h4��J4���Pأ@(�?Ji��L��                     4�D��iH�  @                         z�$B2MRyM���4mOBi�A�5�   z�4h   �   @�    "I@ 10  	�MS�4�4L�L&�4OM  ����@h�� �	�4 h���FffI	~�Dd��n|Ά���¾��oB�ow�}Cនܫ,������Fil��C7d���zg��2X�tݹM7I��>6|�-�ݻ��ؗK��0$݌���,쯭���uCx��v�g�溺�{��7m�����l��1#�Q�͹)%��l�|̦-��׷�ēz�n�m��%�.��A�ώig;l�u~,0=잹�7	�_ri��w����=���v^̈́�<���ϟ$�vntd;�&��[����p*_}c<��{����0��(
*-RP�r�ea��Yki3A3�\�ZLx�"M%����D~q��w�����@����!`#��#}�8|8)�AL#b*�5�`)#�I���G��G�cI].���!|�P6�pT���༔�e �5,�s-uKjjA�S�Z� <4�Q8��$�"
������@@Dr=�P5:�Ȝ�ЈNx��.����'�D��xgit�-E��]�ȥ]$@�Q���1Y��&;�H:�~�,w��B�ۃ�Ã 0�f��4�R�Ij'�'���o�.O��gly��4ͫ�@�����w��<x����W]�o��;v�[=:<����穅�5ݧowk��x�<�k��wz;69���;�@ �(83�,c�%Ko���|��~X��^)��Au�
A
 	U�����4�wە!Ϧ�����Z�Ҿ���G�/.��b-_�����յ7a��:y�<d�hjylI"L��wg�vdؙ�a��P�f	 JKOTu�����0�!@�1�&@�iz:�`�{ I �)����`��I(iCz�T3$�.7�FM��i=����1�G���k���Th�|����Z�)kGM��kwA��_�����||/1fXT�a�$��Ņ�$�4t��������ZE߆fٜ/��&a	���*Jou"[n.�G��E6)4�ֲX��z��A$��cT�D� �kH+�+B��k�lޚT*�l�ª�X��H�U��i*5~��g�K��2��脙������Ӱ��-1%�HqP���]quɊm|.K�Y&ϕ��� ]��P�}G����)X���!�)=������F����!�'����ā�XS�D�I{��	AA��!S�-���!���4���JZl���EbPR	K�ا	$]1gE��a�sQC�f~vr����*�*Q^��C,�o���M6�CG�5a&$M�(h�b�'�R�"<;ݜ��ɧ���c��*��QD�:�RG��B�����t�]�x� �
��Ț���%� �vA!|$m{�w��'�}O���'ݻh�?}���Ƚ6�`CA/ �IG�_c���#��(�M�%�$�Z��FƐ��L�����$')�G�р|:�j6�Is� ���#d�s� @<�����,��3���OW�ު��W\Mq��j[�,��b� q�� �9�Da����r��삍�����������poA�p��0W��ٔ�$�o���]�ǳP��"H���4�>m�&�O'l�IIs�.[�A
�5-���\��7���n��x��w�9��?r��$��Ѣ��Б�v�ߵ�  ��@������?`��$e��~~����]��r�����Hp��K�A��s$Eڷ��	��mKXpQ4�'����_G<�Z��MQpC$��F��a�E����W��ϛ��x�`$��`�<Z>����f�8�Î���?�R�\���B�u ���י�
v��F� n��Pd1���6I�M$ �f~���}w�>��ҽ��w'��8u:&���v����s��T`#�hb�J����-�Vd

�n�S1r��L+��A� I�2رU�t�`���;**��E��:�z�%I�gh��.m�0iKJ(@�W"=���ڣl�@.�����&=�l��~f
:�J��V��7(��RP�@!����~�ݬ/��J��H�~����DN�ʰ��$d@B �3�~�׹�܀L9ɓXi��fgٳ~�0��4pp �F��4
/��%'�����L�3�C3O$>?w��5�Kԓ�<�|�J=���QX��:|����(����Dg����pfRR��8"��@�SUt��yr�!Ό�F�:i�b�B!���7�.eS ���#��ˠ����VH�O&�� �p�к�@QQ�X�`0>~!A��r	��P)��~s��J^6� ���!����!=��i|�q>WW�DYMd6��@�֑m�C?��
����~����)�H�����e2t"O|0���� ����>m��|`��{ĥ��A��H@�Gk'��ύ�e��1��B��҂�T2�݂�YĐF/����U����sr�@�x�o|c���= �|S7�U(�I7� �<Ȕ\�;��b(96�0730�Q�W6�?jȂA�Ut��|b���]�o����_�pC�G�܁7��˸B��H��ɵB�6r�d#uv겍�E)Y���x��e8��.��$V�T�TOŞ���tn��t�OQ��饳S �7N��G۾�Ԁ�c�1|z�:k���>��1�Ct�vKaօu>RF8"ꨑ�)����/1J,�2��76�2cOT�PF�E�7-T��T��(R��,"̉�_&رu�FTLФb10��߾�:��
:�\TO�*=2���Ɋ1�I�* �q�ؘUFZ.�����{8���X�?�ҏO��;��e�|�k�=����|)a�g��(*�/$�,���7G�	�[�6I%�7���:W;)�ӓ���3������{�}�i6P)A/ke���u�ld
s) �hA4�ѕ0Hk�.�s�wRB��C!e �[E2ӏ0�S(r�14�X��a�r�$�&.`<��fM7�!o¾X��cU32�� ��2F2C$���q 3��Yռ����e�X{{�¼��6��D�pp��͂bn\">�<f��o˔�������8 |h���(�jSiÃ-��H������M]\JG­*eiE7��8�@l�w}kI����T��As�ö�Ѓ1N�I�S��:�����$�C�'�2'ob�ښ����T.����,�?u���3��L����E{voȤ�����50'x��l3���]���H��Jnd��3"[�h�/'��U�0�}�f��	�[���;Jf3��|�-�mBfc��c��ʄhz�}�3f�	NHG�L������|ү'�qq��$���7��h��O&�s���Δ|3Q<����/I�����(D��1����\����=���6��E��va�>��	%Đ\s ��%_a��vp�2��3��rR�����"E���89�GY�þ��s	F_�?�����p\w%��YT�gƮ��P'�@��YX9�����q��ώ��xt�ŀvL�:����j��8D$D���n�_?�=F��ϰ�Y�A�!*M(B��i���%� �����_)z Q�#ɰ�� ޡ�n��??�w��@>~��~>P9�j!S���O_��w�bdI@��Uh�ףՋ4��~�S��q���Q�x��iO����w!��l$�r�8�>),�5���T������6�t��L���K����90\�2i���� �����G�K����Ş"�ZL�3U�"Y�4���HC�4x=��<��)�@��2r�� ��@��ҳH��mp����4��ت����&�P |��.i��\�X�"��Ɛ!�������Q�i�71��	�����@��E���֌�&E�����c����O{%�8W������,�[����M�n,�8���Xb�@�N&DIq�1e7-�k;��-�gC�YsX��I,�%�H��s�rD���IA�f� o����IO���q?+����ػ��sv�2ҽ��+7�Yp��Ռ6�7"��ϒ3*E�P���������%�I�I�4�ބ>�ψ,3����w>�>����6P�g�G�@ ����T�@-�~�p�-�w(u��/].�2��Iȋ!G��&� �<��Ik<(�!���x�ST��g���Rg�I������X	!y�U*�c��ŏv��
݁p��R���)�E�k֚��e�����39"Xgء3��@����ˬʘ�JR?"�g�Uf�IQA�A��P�� M�)�"&� C��%E �����_(ԏ�N)���4I@����Ӹ'��Ǻq�17x��x���_iW��"���D:8* ��؈6��v<�ʗeSW8�*H��f�]���?cc�gTɩP�>4-�HB�~g�BhіM���Z��@�FH]�%����fж��	��l-����0���&�wn )H���
�K�W2>ט�.��}r0glaUJKPqyMG����C[XAВH�9ؚr*���i! �.y��S���=��f�>eb�j
��1O��	df�+�'#�ᗧz0>.�"��!�"7u�X�\�oP7�'W2ފ�5�ʑ��	�(���$,!Ֆ.��Tn�Y��n��p�Q��ǯ�=˕����TP8�ѻa�nc[�J��ז��y��[e[��Q�Qv"�/��F����vDWe	��Pf���@���^G7甤�0��A�gǾ�� xvۆ��n��d~�o��}�|�4�.}F�z7�p�l��P�);�R���Iس�Y���$m.�"DS8P�A><�Y��7d6ՄN��X+ad<Ytxh ���������:J��=��0hY��ޘ�N	J��r���(z�Z9�복���+̏O����N#ɑ4'?$��5���C�~X���K�Ɍ�׻��f�1y�6U�m"B]9(ŷ!�[���)Jr*d˘�G���1P��Y�4,9!�v�ֱ�]�>`7�IHn�$]�&M�߶�a�u�)!��η�ҧ&�)s�|��vq��'	�HW�C@���erS�`���"o�f4�ד����"�Љ��r��
,�Q�8�*r��waXā7�v���yt�솨o:=t��[;�R���	hlTyF���b�eAdT����I�oo&FS*/n�:��0�諫��H]!l�s��r�Ar� �����DU�����R��ke�m�-���X��j���u�����R�m�[�kUFƤ�6�Z4U*�IF4Rlmɨ�$Z,d�ҔlY��ƌTĩ-6d���l��F"�Q��*=�!��m�m�Ŋ���۸�E$B�����h�(�!��L����E��#�$�",`���T�_d�DIAv͎矎��楐q�A	ddTA�Y�GeP"��H*#`�E��E�$ ��R* �@B*�"��W+f�<�%�re�p ��?G�l���4:�M���Wv�{l��?I��k�� �ٙy��<ɵe#@�dAK�d�l��̅�]���f�A"���b�b,��"E$Q��E� &��b��ųr:\�@m���л�0�ۛz;�m��z��߰�ƀ8{R������������� �ٚl�-[2�>��W��U�D�>Ϣ��Y����>U�u��_����},�?nc���}ͱ���=9��̿��?��W�{�������o��?V(�"}7��R�M������_����q������~w�?��i���?�q�ُ�������~�O�#��?�}�����!)=W���'��/��c��С������-��Ļ��>��w�nX�,�����~��ߓ����
!��G����L�����Gy[��:{��?������%L��=W�]�2?��t}V�}�����61^��z߃�����K�M�Q�g��A�?�җ�>�����������~w��?�2��x-J����_�O��M���z�^��p�1�{�qZ�?|P�J��T� ��m�W�8^X�� �����w]�}����#�>8��o�w���o�Yx�������y���-�/wO>�C�?��){J}'��>��������{�Gg�~��W��"�)�|�u)��	��|s����iد_�^���n���}��������X�W|?q����
����~����X'�,}���O��[X����8ڿ
E}$��}��C�����s/��~K|	����e������G�}/ѻ�>��g�=�����C�כ��G����C����_������O�@�K?�O��6����������M7��g���>�ӕ��_״��,��|Μ�=O9�a���{����g���t�W����2O�o���8a��]�cI�u��&��f�:�������`Ѐ�P`AU����PC;?W��Fi����۷��֎\�2   /k�r�L�m'���� ZO�jJ�to�&S�`�sx�o�O�+�f�O�v�ps�@�e/���8�����bdQ$�V�-�g����i8�p��M�S��i����aG�4�����DJ�ާ��pw �6��&:89��v�Mm�>޲���j|`#��ݚ\7�|��� �w�a5嗶���t��9��.s����J�C�����v�i�����2�[��Lzy�&��y�n�C���D��΁�c1π pp�|��2]�8�_'�[�#�]>��>����9�ZR���>ߕ5A�0 s��򽺽7�>�P �t���x�úƙ�z�����d�b�P�2���ߢv���poκ\���{|���k��O��ʓ��~Yk��e�޲���e/<g��i�^0��W��sd �	���C���	������o���~�~�^+��[���΃�cM�A�U)�����K���b ���,F_��{wg��O�2W�ËV�S�ܿ����˗��}h���L�C1���9���8��G��2�>|`+�������%��[��+��}Q��١�Ә�\{=����}\��2�\��/H.G<�4�M~�hɿ-Z��Ε!�V>��s��Q�w{�}�ͷ�{�x��	t��Ϯ���秇an��]4a?��)����E���W���gдIg�m���t�3���)c�ƙSI�ߧ�� ��Na@�?��?���v����o����vQw����>zJ9�������x��vR}#ƽo/��Ѯ���m(�U���pw�@|��6��M=��~89� ds�+����p�b������'I�y�z�BM�����{��딹ppp��(H}��B6h��޾�v���:�0<��c�N�D�Uӭ`�/�>>�U�H�9��@�b� ڽ%� �1_����G����W�JK���v{������7��^��}�k_��	�#F�Z1��6OXD-8�_�[.[S뿞?�����u��8��C��6�V#���jtX@?94z�u�s�-h�N+5	XVƩ
�MR��^�Z�,t��k��v��p 9������|WDχ���;z.��~�vA�xWl��}eظ ~6�Ͽ��ۇ�Q���V��{���~���������F�ʢ��h���!���$���soiŊ0�M�A�F��>������ǅ��M�����88c^=�������-I�ii��Bu���s�e��qu����쳒}���Gpv��8�)��vټ/4�4�F�ʐo��z��韎�v2�r?�׷g�~җ��۠p���T��1������֩,��<w 9�i���v�o|���!���e�����_  �8z��~���N�!s�������a��龶h;���g�l��,iMz1/�~�;W:�K.]����W��Q�X�����!���w�(�?Ɣ�tL�K���8/�l���Nݿ<��>x�W(��I����?��[2*� 89�x叧�����^4��-��z��hpv�9��i�g>o�y�),S�{c���s����y�/�}@pn+�Κk��u���o��*��~k�sF�Yq��*RS�����~z��!��8z?��K<����=���zۧX�`M�O�npt�����p�������a\�9��,�/��S��M��=���n!Ʊ	����o�硕��ӯe���j��l���?o�@�p�|~��x:c�����mW�vg��~�k4f�;W��)�6�m�r(h�M�XZ*���QdI�s�����z��0�-*�\_!�� ��ޡ�Œ>�g���4�,�pǴ�:�i	����ϟϦ�������N��+�F�|�Ӟ}�N������c�)����ΰxM��������ppp��+������c���{#����5��Dw��h���j�s��p�ʊ��e�z��o���"v\{�4��_K�9��݄a_�!����s��8[�������*;�#��D��&�W�ӻ���^�����/W9�����'?o� Aq �\p!ie��ъ���x�[ڒ��~�p K��l�����ZcD����_Šl�⛉$O�
��oπ� �	��g%�Yg��p�Q�4����������M���z����89�O1K��q�gi��m�'��z�`��x����Lџ�geTﯫ��I^��4����a�89� SLS�׎��=k�Ea�m��`ۘ�d���o��v�w�W�>������+���Oyk�qU�j�Bj��9��-�*�?V���\?�,�Q�o��v������ݿ>@w�9��O۫T���8�G�"t���B�hv�/�e�΁S���������88v��{���/VK�l"E7�Y��}���	��Z�Ӯ#�r�j��#���=\����e?^>��kƒ�l89�!�����c<$-�lܘ��z/��+�Բ����p�-]U�fi�濧����8�888O $���O��.^V��*�o�Jq^n��o�>�ӏ?����� s�ጸ�s��+�����%l�`��e�T�+5���~�Γ���1|��^߉�~� /em=����,�/U鎽+l��;Z+�y<6�����R����/���.s���Nlm�-��.��E5��`�����D��p^~�a��	z�������z �8Jт�pE�;�eEK�U�N�u�u\�4�话AM�CR�9�v!���-������z��fb4��:K7�E�J������=�| . 8br<r��ja~6��L���G���
wO�u��I������Oϣ��J74�-��e�{�	R)~�P��`��)E}�}?:WJ��XB��Às��*u�|>���)ߴ2&UX��G89{�L���l�FO��W0+2��T0��s锥>��� s�!�iP�Ɯ+��CmZ�g�����s���������(��b��k�v�6���tz�'�P��z9����b������|sw�s��e�����n~����rj���徟���s���dr#�-������u�,?/�ߴ3�v{�e�z������a���3��I$���ѧ�L�h;��i�/3]4ۍ�JL61R<D����.orl OfH��`�f��O!�2��:¡��V�D�ri�!M�3����|gv�J��zROs�-��m���-���鸲��ɭ�DѾ��t���d�F3Vi&�4�,�]`�aac�i��Eޛ��'N���8��=!8�!=Xf6���ѱ2!,}�t�	�Im��35�y��T=�۽�9�Ҷ-����A�:\n;�E�Ŏzڒu��"Dͮ`�,�e�f�,7wC`fS���ǘ�\�nI��Ҟܥ�ǰ`U�n�JJ��wC���`B�M��j�������.�m=f'��ɔݛ`%�%',�D���J0öT�5�!�+'n��u@�X�����⸠�P1�qnW�Z]�'S�IM+��ĕ��B�aN�\Մ&�R�H@H^�` I+���xOO��W))� �Gll$!�wZ�!�ݻ5p;v�n�HW�uC���!��f�e	�WLǜ���W O)@�Q4�tBE�m��� �"�{����R�H�F��r��8�b@����C�*9�x�B+:�C�M�m��y�Xɫy��-j�՜i]h��՚l��e�����$��I`�4@X��Z�bVi4�Y���+�Ő��В�k�(�n:�m�Bh(D��vn�T�]i�n�d��m)9i{l�b�%�K	�Ag;Jӄ۽w:ù�ii3k��T`!�Q�V/6�2��YN%4d�,��ŉ�`��M�i;,xB�fƵ�;f�b@���B7G.��M��z���6��Ê����M	�l�i���c�����FX���� M�Yu�ƙT�F��v݌A!�4��!�X�Fu�Q��Sl�7!A�M!T��B�Ɔi�˻��l֍6Ǉr $�6k���t��2�$Zz�Yk��c;R�v�a��pEH2��R�4tk�m��i+9����Lun���0Հn�����p�B�Hd��e�F�n�%!��\��9����c���IB��B���Iwe�`L�a�Y��^��e�P#5�k��z��l ,/mu,�I '�^Y:+�ɦ���j�s��UHIČ#k���i;dq8�)ūV��{�I�ݴ�'W���5�j���ffwM=c ]�Ѐ��i1��e�e)�S�,Zn��IR� =
r���YI�[8��5���$�1c���aH�3l`
��q�h�x�@�q@TJ�p�[���a9\�D]�sA٩���{����OzuS����ua%f��d��v3��B����\��;��є�!z�%����rz�t�"D$')*�Y\rj�m�
�K�v��[.X;��K��WE��V�&n�#m����b���n�&�W��5�Yx��)M3nl��绎A��q�t`a�CH�1�#�bGFy`=n�Rћ,M�+�8w�;mU�\�ڛ��^�ac�q)2��hD��F�n�V�@��wY܆��u�*Wvi�C�b�9�`��
�>W��u�7�'^�(ȁ�C�'R���� 0$*���&�L��撮���i���i��77+AYH��e�����X�`ͻt�,��t�y�@F��a��:��y�R��A��n���!	b���7���JN����,�us}2�u# ���KY���6��4@��%k%��RZ��{Xjg=�{�ڝz�B��5�N��X��qC��W���l�I�O�3Ї���h>I�5��E_d�M�����&M�o&�I^�$�.�*��fE���E��e?�I&d�L�$��۟%V�zL��S�N�>�ﶶ�mFն���3$�,��$�~�*6�k4��!]�k�$�@�M'^2�qs�1����l	������u�5eM��e��c''/,������] R'�̠h[hNZ�����eq1`BcYݳ����0Z2���lt�ڶ9g�g�AE�$�{XJ�gk3C��Mù!�a��dLt�@��ݏH7{�% �@��ӊ$*H�a�B�v�c}glNcX�Ƿ��L�`i�	��k�����Y�H@��|M.�������Px��i�M�%�ړ
Ƴ��0��Sk�{�iM���sz�w��
���@�+r�u�b&�  2C
��X�Mc�ˤg�Xy���¸�I)�𛦙@��u�)$I8�	��\Q��/ɸ��Ҝom�+I�.���]���62�4�A�8="����o�P
�'_iC8Id�`��)
��f!��,M���)p����ϩ��∳�BD	&�,��Ї{v��!U�q�����I�ĳ��)tv2�"ޜv�ri D��(�F<�U��17w���;t���ps��؈�.)eI�$�V:�����a��ku��];��eέ�$U�� �N�`H�N��s��	�1�P1�D�,@�i(MP6ù�!��{�����u�z�N(j��0��%�.���g:gA�g�eU�x��54�C6*��;eݲ���1IS�5]�G����S��C��x�gg��X᜞��ID�e�(A����x��'Bajo%��`*7#���,�J����JF�Z�Z���E��"���W�f뮴����0�$��Z	Df�8�j�M;]�����Xłn�oYH�]w�޷�Q[�`B�`mꇣ<M&�\���s*O=Hi�� �)b b������CIOk5��D� c9e%c6^��RZ��Z�erҴ�[`I�onD�X��hM2wM���B�\p�ɥ,���ji��6�'9k+	�3��i0��kT�6�k���\]��Lv1(�Q�\���Q,��r��'�y� EC�Cv�Yc�-�����H���%���ݼ[6Ft��ei^�ӈ���X���B�ۦ&Rņ�K	��wr^c�P�����2Y�2�UkM;��fք0��%!��yЕOt�ij��7�vUv��K��a���+)�偬�mG7�%��&����싋�hP�b�)�\5Hx���m�v��-b"��15��B�Z�t�v�́V$��6���\�@�F^��Hы�4�� a��ݎ�Ŝ�V=�% Lp�K9
�1��]Yv5H��,�'=]6�$�o7Y�`�wr�]]+�\�r��ݳ�k�Gkkե&��s4�8��Ec�L1[�ښbJ�+���kݲW�<$�k�n�JK	�.�q۶[�en���R��UT@1e�!	X� 	7��@���B���c��ٞ2�Ha!6��  eq�wl*mYL�Ғ�SL��@�
ɤ��s�7Z��#�0�����B ��e���s�h@ �,�N3�n�oe�8Q�4]��<x����Mc ����u�%$�m�ݷ$�m`�`$zY�B�g�/֚�$v�Y�Hk��Jp�s���w]�u��p�ᚻ�κK��+K���s3�r��V��e%�%���@0!9�3�3e[�� ���3KG�,R ��v����#�UA6��Z� �L�uhZ�QgZ�,�	H��V��Id�����C��s�쭎Qq�0� 5Mv۔�RJ�(Im�٭��U`��Y�����@L�"�m	Ad9�
+�nD)�RJ�"��wb�"T�+� +�
�"F�WH�՚G\离�"Ki�e�@ � �;�	��n�CV`�ZE��T).R,S����¹0��6� �X�"S6��(rYe#o;+�Z\1�& n��f��8�J���vF�."ac8d	LV$� ��2��S��6$�`u���DѦƅ/6q�$��6lB��Jf��ݲ�󓛑�e�x�F "��9��wZ��ݸbb�G4�\Җ�A����4u��c��x�ݫ���� '0ֆ�n9Qj\H*޽��3p��L�I�r��2���1	�T�&NjYb�BRB3��bG��l�4!4Lc,D��i���KH��fĴ� %0m�AD��b-s��X�e(@�[A��U�6�F�"XC�F
�R1&��9p=�S_��U0 ��V K5�[�U&8t7R�췘�HA� ��+T�+YH��ZWY6���D݂�e����+�%$�YM0*�k:�У�X,&��c��2iM�I�U@�S*�Zc9��Y��`
[D����3�%;�9I�[�ݤ� �v�&�Ơ����{��a$3`�5�CX�p0��X;r��Nf�JD��0�3-a&$+ag[HW\f�IT�ͱ%�M�������a����9���x�sf�+6�`���II`�^�m�Bb�+ʰ��ٺ$a[r�\^��g@�Q�掛�Nan�6�mR$h3A��n3X�)�m1�&��\b���"����RKN%9��W�m\N�!M����vɫ�W!H����i/Ĳ�Yzwi�sK	�IDH�-B,z�+4��M���q�����f�����lAU�Bp�Xq�+l@���=vYâj��C\�i�l��2(=��qz�(��%'jVim���#�l�I�oooT��/VJAX0�sl�4�]2���P1�,�"��U'wn�s�JĈ�D/=e���=�]i6Vi�(�����"6Ԋāb����(����c��V#aK�ec0%R����e��)�!	T�^��$'�ݺ�-��G%��a+��Cń���v\�u���X�^h���uf������40�Khws�����Hm�[638`f�"`��P���GV�Kq�%A�X��B��,�ڵ�c�|� !��Z�l�,�2����Iq��*�R$�-�,Y^%P1F��i:�Mv� B����'	�z��+հ�-
���h����v� Fk���i��Q�0� �P4]w\�!����^w\h�e�rl��:Đ� ��(����ji���6�u`��1#w�4�M.��D�[J�f�J��] =���9�wXsK�@�R�Ts0Y�)#��m4�;��x�˺S�H���Xn�p�H�� ���D�w��C{]�CmY��P!�����{d���n�2�2L����^���5����޷h��e� #Uj�۶�)���D:���X35p�8�M�<�{�vkꗔ�3@��v�b͛��h ��D��sx��􍾶Ε�f$р�]�$_X���J���D�İ1�{S
����8! C��yf��urJ���pb`H��!F1��f�*�3�9�Y�	��	�t&%\B���K))wn�-"b��	55�t���5�E���%(Vo��@𾷡���8��x�%�7@X�@�7}����c��o�CL��!C8����[a`a�y�9�`��0'6[TtӍ	�6Q	İ��B�Lx��3L�=�SH� k�7I�Ge��⁄�К�d�۱d��l a�r��B�oW���fd��(B�,Q*
 �c�
*�A�,�"�!���^,��&���kJ5sV�}��/�7[��r��r4s������wv����y�r��2\�-r�����.��9�D��r�H��X�w[�\w&�r5;�+��4��&��2L�v3%�[s��
W�)1$��Q��fΡ��ΌG7.��]�W;�H�DH�2"ȑH #"��B����es����x˸5�my��~���J��_�;�}/������ݡ�ޯ�������%F!i5[��^Q�c��L�tߜ*������D!"�ͷ7l���n�h۵�-����eek����F�l�dүEI�YńSG�ٓ���g����"fFs³��~��EcE$�R�|���!�ٿW���K��y ^@����yy "�NG��8뇚"@`�	X�e8�  a�� \�����-0��s?�;A#�ߪ��|�:b�䭢U���[�[�	��c�;r���$3U����C�9(Q��G�Z|����tOTTh��=�``Y��|E�D	�ױ�}�|��Ler3�����G�G�P��eh$�8��$��&�X)�,9�<�`R�<�0'�ԑ����9QL&��AX,��{���K��1��\y���k��{C���\�_��+�� X����'F��#Q��`�pԅI���
��WE�M#��>t�sZ�]��b޾��!M=(����ZG,���
���(J��XW]9�-�`�p6�'2�v�`G�q���}V]*��HՍ��%,���A�2�먺��>ا�+����c�|�8m��F1x�I4~AmT�i��6�	�Y��-UU\S�J��NK�dՍ�O���o�N����w(�^ zQӛw92�<�Mw�	�[��,Cd +K(M�3�&�z<i�&�<!�37ygn^Mr��ϱV�BOH����>���|�Ķ[�U�#�#�L'~8�Y|&m�]��z�F$��q2ᔡ<NqG_N��P��y��*�_</� +�G����g�(;`�H���z-D4f���E��C�D�B\���0�9K�J���1B'��� �r8f�R���*��Q��,��)��?�"A1��Q3̖H�U��TQ06���" ä��k����h��|3l�����TB�kH�q<�j5/x�L�9��b��nH�kt�����uCJ�`c�cI�:�l��� H)�EE� ŗF�W�勳!�,V$"������6r�'�^�!�>*��)35B�f��$��F.1$�`���F�W�:���zU�P��D0�V\	m�݅HR��Fȫ1QΪ���]mg��p!9(�n{L�D\<a����Տ
��~�k	�E�FCΒ6L90$&k�[�$�9�P�dR������뢥��I5��b�2�XƊ!^Ep��T,�l��� (kr.D�,��r"�y�K��;T�n��m�)6ࠫ���������,,�#{6��6m��ү �8QP$U�mo����H`�1I��bk0#L��6DFDݭ��(���~yU{m�h)⢊!ea�+���
qT"+�� �U aeX�a-�幾��������?�i^�ڤ!#! �D�L0AA(����	B�b$Y!C����7]�>W��z|��ɹu������:l��Õ�9�Z������}��~�F{TG0� ?�~���뿻��U��'ݾ_��֝D*B�'�1>��Ċ@k�O��	M�wT1��D�	���@ ������>�r���HC��Г��c�k6[O���"���B�o��bf���Տ���$	l��L����X>k����8�|T�%9��d�2A���<������%@s"�@�hz&����~�����L���wWY ���|X�2#$.�����f0
sĠ�Z��,%�]��.%@^ҷǤ�,�F^�(IG3:��Hj%�n�9:�P�3@l�#X#�RԘP}K5J�5�g��Ru���f_c{q�8E���ZJ0!B0��a5���
ښ��A��$�)�(
<4�T5$x͛8T�G��
��Uۙ�vYn2�Zt���`�U[%%T�9]7�!{\�e4���x7��_}��A��Eè
��;���gxC'Xn������_[�Q����ɳ�qJ6�Η��d��e��H;`)M��f"�Д����C�HD��d���3��-�!D{�����9�.�ܕ%w�.�I���ձ������E��ۨ�:OXb1t��%�p��N;���r�s��!|��@=]y��Ҳ���QR�+�O�_WN��7��m�&O�S�jL�Q�X�h'c�Hs��"��L!F��O��ۘ�~�=����'+ۦ��=Y(�Y0�,ǂ��8�5Ѐ�"2������P��#2��]X�S�Ex������.EE+�-��I;&�m��a��m�=�@��#� @�I�リ��iF(7RM��^Dy��$�<q��#�S���j�_9 9��ن�2��������;�����c���PLncٖ� �b��+h`i�1ؒ�7�@G�D�GC�*���݉H~]�UC���a�nQST(��);�����ڍ�e�ë&ԁEs/�I�]/!��w�C���2|��^o�X|IE�3��V����X�o� �n$hdYr�l��y+�u 1A6="bE�*D�)��Ա���J�,E�/(�rbUЄ^���Sq���bc��*8�Q�m5�	ѱ�K���«�0�q>�;b�˽�:���Q3��]ú`��h����á�D�����j�I�����m&q�Q��(���WC��yB���O)��aħ���S�.�zZɊYS�s��g7�**JC{��\���;TV#�*��[�|e��&:�X�G�Uxܤ�\L}�UfhL<w	#͍"��kazI	�����X��i\�Ѥ{�;�ć�NZ)��0�ko6�Z�g�9`�!0�
n�qY�+>�G<�I:YM�nt-Lal	2�n��F�=ה�8"B��K�㐺�ᐛI��Ny����"1��<�0�S<Hh�=��v��L�F3� ��M��5R
��T��ND1'�5)2³G�\<f�'�g�bł���N�~
9�LW�hf�H�pe>4\��$�	yK��Ԏ��ZD;���6L��qQV�� ��4�:��Q�u�����J����,.]	T���1åC��Y v�δ!�y����"	���[+&Fzx�<��ٱ��dO r��3�)�2e��I�����s�RG�0�129��%@CL�E		�^ 	F5ETb.��ҭ�~������ot��|����Y���S~[�Z5�6卨�9��h�Z�ˑ\��X���*�z+���J�BտZmkWM���i�U�ԡ�#U�E[ZJ������t����-mk����}�W�6-�KmZi�Q\ۚ�*��-�7
���m^Y}�sW�k[\-�UҶ"�( H ��$`��-�8%M"�9�6 �CP����pD���H� ���(�b� Rb_��t�h��(�*�R�	�ϑ��Q�ѯ�k��5��Z��[��5x�zU��4uATPT�.���n��B�����
H*��T���O
m"]`(�!u�Q��a� c��D]6��f4��}�o�[�W�#2*�ԑ$t�c@���!� ����"Q
" Q(�@�0$M/��Q.�����*���SIc4C�4�����k��A���^���?�d��#WH�G��߫&|��X "g��QWV"�Թ�P��i��W���-�]��3�k�[H��M�t2�����?/��.�Q�:��D�kU��;~�Ť�Y���B����e� Ȩz�~3�l�oM}�S?2l7e����C�v/CJh���������͆��w߭�,Jg�+��L�y�Pu_U���D��,�_�s����H@ߢ�T(�ȷ�K .]�@R�$_�绚���Vǻ��hd���@w�;j�#~���+��eh(�:�AA
ET�@E@z��J�NxX+�_�cP�h��{�jh�]�  ��M���㴡u�!�y�I�ki���y��H�o��S�e�{s�r��/tδ˼0�i��������Q�w��;;|�6o�?�����9����� 
�r��CC���M��m?�oٷ��2��=������n�݇��'j5P$Y��*�gꆧp�����y�CS��ٲ��n��SA^a��_���&�u����=9v����s�?/������{���BL,hn��k���J��eI$PE$D� r�EA�D�0U���x�uPm`V��)u@�P�\��D\U;C�
~d C�� ډ�".j���]Y3UUz���S͚1tl8̷�.AD�8A�j a��"g�M��r�qD�)i�j6���ҕIl}�;�%YRD`Dd	F$���44z&1A�6�mt��vb�&؂߀m��؛^��߻��͵m�KfZ�1���uk�5�cmZY��RlV#��Kc��´�|��mr�ɨ�*l�֫&�Tl�Ǟ���$Z�%��j� ��JQkҹ�Y1cZՕ�V��Mlj���S-��ڻ۷#=uZ��oes32�2�f���h�̵,��mX�֋�5d��ScZ�WM�V�e�ֽ�rֶ��2��-��fj�j�4Z����i�ȭ�=�h��lj�A���Z�[j�W�WCFɬF�������W��<Ut�|\���4�Yx�F��Z-no����Փe6ƍ��JմE2V�Z0K�T�Kb����B�5��Fֶ�5L��Tk[Ej�5	%F�EU�^�疉�nW6�������i$֓$���m�]WY
� AU��!����(E$��Fֶ��Y�+��1�R�
AH]}%�.��*1��$���@mF��Ej����TZ"A 1y���-H+ �b�PE�,�7��woP�����ۧM<[7މa
OV���� 2�ۺM��T202#��2RCEyK�,���Y�b_Iv3�3.�$4-��	d�d���Ō�'љ�Z+V6صEjɭlmF�������kj�[⵹U��ִmV׺��e���"8�T@�*T/� �Zh�fII�38�$�I!��k�$D,kQV���m�m��ժ�%2I �H���8ɓ8̙�v����{y+<{ф�-��Ǯ�����e�U��S�㲧���͚����r�1o[L�\�A�aݴ!5Q]%�����WՀ�^"��p�R(�_���@] #]'�͕�c|�ݧ����z��t�gV����a,X�]
Oy��Zٷۏ�Ҹ*C͗�/Bn���u�̶0�.��
�[S_\k7*j���r5��M&:�`��ғL`Ha8�m�@�0��Xԭ E�os`r���팃֞�MӞ,+�B��{Mk�p�m��l�����HAm��,]&�)'6q	�E�Ӷ������ʰbf��Ҷ0��hxAݰ��Ngu]����>t� �&)�9斏>����\%��σ"HT	�l�a��#����+��'S:�����t��<�#��W�z�6����G��l0�:Z� !��fCs{d�o��x�ʳ���Z#��<@�'���X@� �	$�Y[=��=�J��U�$PW$'�t�2&�J�ubN�Q�
�"7�6or͚j�V'�C�<��D��UO3N$�B:ӉN(h�h����+��;��� �%pӳ��5lV&J�����P�&6�GÛ L"�S۵�G`�6ᤶk�e;�Xf�/�BMQ����M��l���i±�a�f�%63lٻ�����:ʘTm�Be)�J�e@��VKm�BA�R2h�S�����@�'����0������|n�!:$��2�k�kL�>Z�$Kχ�B�V�u�Rx���KZ���{��z�&�p1!�Yм�,ăA�H�!��3��˳ӓ|nǎ���y�$����\��\
�t�0$���;����k��s�M8�c	d!��m��i4�Ė�'�v���x�	�v7v��]��vٻn!&���3a}�Ն�l-r�=ww�a��(�[��<P��4�&�՞bu�����;Vܕ�����"�T�ħ@��m�=�XN1��o]��aI��9�鷃v�ƒ�)4�M���bA��=��x��Ā"Nh�M.�x�R�7\F�+�m�<�B.�{F��o��ࢌ=M�v9�[��p+����"Xuw`(��WV7a6�dL��ye�bj\��4�����|�͆h���c|Kw��i����؜�̗YW_s��[�۱3n!b��uc��4*��LDïn�`:�#	� �v۰��J�B�n�R���͔����b}z�0�wZW�ʄ飔>8�̤'���ӂ #�����nBw��8�U�a9ҙL�7Y�x��=c�o)�n�:C�ě� �, ��t��`\�I*���[���*x}�Y`�k,%x��ye�͆^e��a��*�����L����u�e�`�
��8@0�k��Y�D�|GZV��gO㸞'�-�&ńH�4�@!y���I�1t��r���]m�\k �>)���%YaL�۞'����b,��J������TuBJ�J'���ٮ2�[ �{l�+Q�*ÙaN�XI��.��ľ�䫖 Bil�fDw̖�}�<M�䍲�څ4Ā7ZIF�y� ���7R�j�ZE�K\<�F��Hm�HB�,��0e�{����7̎�l�ٺ[��bi8��h�n�� ���bK(�3�鳝�+n�Os	ʸ�1@tw[k��_I9F���&�g��P�B��S8�V؅�);X;�B��.tb���B]�k�&�-$w[����o �����ŏ���7�%�p�5�u�	R b]q7<N��_j@6�>�&i�B�1N�f�!q�^�}�N�kz��x�x�r��g��i�����	9��t��x��j�/!��lqc�� M�Ľ�����)��4�۳b/�Ba,��vx��HT�b��I�^�k6�7�.i!��6:	�՘Z�x�X���u�y�Δ^���Eѕp��h�g��ى���f&I������E����\�*�^-W�h�W+��m�x��F�ͫ�r��5׍��*��v�5�0j	|E��QV�|�|���K�ۭ����ޖ���׋{5�:mx۽��|6"�/�8D�&(�L"�.��@	��@"��*b�A��-Lg	�O���#�$�j�%�i=A��]t.�Ռ�r�-,e
�f���F�
5�W��j�6���wu����Z������]�m��b��5*�k�r��Z(���W-�}�'����6���m��˛tH�5e�%Q.tX����"6-��i��b+�F��Q��mb��1��,�X���Z��ڿ 9�'�N#�=��m��{�|��/��̀_�-�{������z:ߡ]ΫYCG$J���yo��_A߿g��O��6��>ga��T8�o~ol�_�8���z����G}�?�޾��_q��?O~�+�Q��TW����Ǫ�����(f{�A�
P��D�.�\ܺ ��^������~��ƅ>��D�����TC�'9ݸ��5������������K��9G3����ߩ�n�\L�f��ۆ������O�D��o�^�/��R����!ݘG�~�oۿ��q����W�g9��!����-ӽ�9.V�Rns�H������<�˜�N���D~�����O�����y�nr��}����*{fӾu���`�Sm��v];��U���5�P�xD;�y�[����#ݗ�����dg<�k����oԿ������=z�����4��j��Rk)�`Cmy����=e����Me�<h��D����C�$gn�Gۧ�������.�ߪ:p��<\$������K%k;Y���C����R^2��O�O+ChG�	����m����~���W��o琯�N^�Q�zs������O�%��mۉ~i�����Z���?~���,�h�s�Z��ra�s�w˿g�1�<�K���M���O-�N|��ۯӈ�F����?��!ĀK�p���~�ů���!�/�\��_�~?W߽����DЖ�ffW0�& �D�YVE@w,���"Ij�YM�Z�QmQ������"��QU��2() "�QE�����8�c�HJ������E���1�L$A$"s��6t	��Ap#^j�vs��>�|�}�����k�"���焉B8��� ��(	D�N���t�$"�QЇ=��7][^��B$c�n����dd&����$#	#R�-�m����D�/�n�]$`@u���		�t)QKSJ��IX�@�7�o�dr@*TR�ˍ������e����
���&)�f��w#�����}yb���1Q%wv���w�E6]z�^N�Ю�O=}/[����p��2���߂�	@�¨��$Y檀$~��d~Ʒ��So��j�cr������wE��@Mp��)ݾ������x�wII(%��� �;��� ɂM�ڷ��^M��b�m��sm�V�-_[����U�m��u�h��]wnS�qݫ�9{�ʼ���w\Cί<��ܱ��d�ݰ
h��O�"Np���c\���5rcmxܪ6��U|Vڍ��;F���W�{�+�%ݺ�ArM"E�>�e d��\I>��x��wL__��]����/�\��R�w+��fk�t��w��7s$b&]n�jƯ�\�U�ش��W(V�n�tj8B��-/�K����x�]ۍ���k��n'���ב�'����CӉ�E�#��u��!wu%wGAp��ܵ���_�?����?	�/��OK��6��0o����_��>G�?�!��0t�>��U���!���/ �������g��{��ž������?��j�����%�߂"���G1B �A���X�ccko�+!�)t�
����n�Q	���$�Ź����y��z�x�#I�Ҋ$�bbR;��^y�s�t[��!��On�^��(ߎ�mj�T�Z�T
���{a��m���.�vf��߳��ev{'��6N�G܊/��Tw}�=�}ջ���L���7g��㜹󯳎�$�3˻�aV����,[�˽5��=��A�0FW��b ��� ��6�O��k�կ��n��p(�Qb��w=;J�����3�}�x���K�%�y�����
<\��۹I�������w�⽛z��m�o:1�6+�9��֢��[�m^�Ux���61X�r�x��,~��h�I�^�$�D���!���˷��z����+�Kҫཕ�,;����i3OS~���̯��{��]�������%V��y�rs�����U_�>O1y�C�U:��B[k�r���z`�F��9�uE���|qw����F�|���Q�%�n�>�0���!ɸ}���x|}]��K�U��B�a��&��$]/��x����r|G52�^ ��3�86ᢲh;��R��I6s� �K//Sd��K������xQn5f�>�p㙇�l����c�dr��ǪŁLQf��Șp�𯎜&�9U�s&p�9�In��Ñ�.��Hs�I�S=��h԰]\A%��L j�t_�nT�~���yƾ��-=��}yQ�g��(Cp����P�&JA��װ�Q���$a��<ˇP�)g_>+l�~�s�Ȗ�BX��ξX[�,�S�s�S1�Q7����th��®r=U/�v��p
bQ�d=�&�c8�v� �S�&3����I+�&c�Ξ7�h]��]�$�Nbv
��l���*��X�Epk��<e��J�¥�okr)���:���	s\9o��]��;fx��q�9{k��L��t ��|��8�����=P,����I�N�2����ִ�O�QA%�̘�iKG�Wī�&�/�d���(N]�y�Ir��[�FIX[yY<�����Jam�ٕ-�"�ϔl��xp
�3�J�h�@��[��F@: ]d#96��T���鰑�l��A����V��ݝ,\՞���$G�$����ApG{�%��3o2I�n���!2
lP~��@�����6�fl-*�PQYN�H���`���Z�<Xe����!B��Ԕ�=����Y����At���ď0u��P� Ӣ�PU�����Tz��À�آ����t;�-څ�_E:�����J��,��U�;$W/ ��3�]��b��㠆󫓒t�������hr$�
�R��d�⃦]��h�N�V�ǉ�!^�+�W�g"c�HDq2}yg6Wu�:�%��i�'����<�����jybBnb��Snq��B#r	��^^]A�kHL:�r�$�n"܈�����ǪzC������yZO��pVt̔�آ�n�H�f�'j�+�N��˼�j?e(�Vys2��c�s�-K�>J���P�Q�nR&xm®4�U��ݱ��ΠN�Sc�A�/Q��g�5�7Q�2jǃ�	0�u��_��#@:�6�
��_ĳ�^�Xd���7�u(|���ˡX��;�2�޶��\�.��Q�6a�^����S�KY7���{�)帼1 ��q��'o�$4���@�nD�K, ��˩����B���΄��>� �0�P�+,\�c��S5+�Y��&ky�	.��������Z�jXpq�qF�ư��A�7�K?G�Y��r�	� �"��LPj�8�N+�|��_��>)�X@Ź���/7u��~y�wt���u�Wo]pR���B����I����[��ŵ�͹��ܴm��m�j��կ/����G�����̑�|=w�%��t���&��Jr�M1\���|�Ģ���<�%����(ƣl��m�b���s\4o�Z��Z��o	���:�HQ��$��뫜�מ\g��#1#���]��(�!)|/<޽s��x�^��4x�;���c��b��*�4|o��lTTb�k_B��涽�}���c=ut4�R��d��w#$X#K�<]F�l��ɞqN�}iPa<#P�a�)d�^���z��r��!��!4(R��ҙ�����wR=�L�E�p�$���TE�v��M�H��;���`���Q�^.b��Z���4[k�^�Z�5�k{�t�{�W�F.\F�9q��v�2/:豾P�W)��^��η"1�����k��~��='��ߡ��O��w9Xz6����_�>����F~�&����7��_�h��A�T!��3 ���h�Fe�_����n5#�Xr�������sH=g��1��������N5 o�p(� ���KP切���S=���v��
�"�<%����A�;(J�ʥL�1�BƂ��ĸKhw��`K2��������!�"8����o�2l��T�l٥^�E���11P2
�g��Q��EXh�N\�/)h���HQ8�����`�%���h����ӺR��H��M\6���k�$o�'h\�������߽��jy�8E)E'��BἭ�&-խ|��*+{uo�vp!Q�`�.�)"��>{���o;,L3���?v��Bٶ�d������щx���NZ6�(i��M�SRT�4�A�h��޻q���2^�<�r`���2z��)��9 +�a�]��&O�r�mM���GL��	u�Ma���w4ij0 �Dj���܉yx���0FMS�|��;zм�GA���I�W�����B�E��ʯxr�gj�Zʥ�B���q6�F��s�	�_���mgtq�fA���<H5�w.�&`Wz\A�]R+([��+�T�xs#��3�It�-�va`b�\+�C�~F���36f�'Er�ت�)�"݄r��l�`�#�F � `yq�@M��	N��(WA��FvƤ�Zމ�C'��fp�΀��R<���)"!pw�i;3ө)+�T�10���Y#�a��@�M]��n�	���Z("� ����78��S/:p!�2�O|
&��VDA)�j�ܔ!��|�l�ZgKߣ]�J[����SD���1NP�11ڈ��v/<�4��>ua�"�sAgU�/�q��r���%�2�J�JU��(��Q�N��o�xS�����:c����x�D��Jg�9*qx��(HY^IWsz�iđ����}�>���^Y�p��C�y�b͊�k3q�:�B�cI�EP�o�c�L#�Tc�QNu)a$��V�?�n��v�*�����o���_��O�;wq v )p@\�)qb-��[��rѭh�T�"
�H�"���  k��+�A�Q�6bn��	$��EI>]��L��)���݀0�1�Q�W�ڼl�j�гm�h�ս������II�A��~�Ȧ C!4���,�E��
�I��#?����[��ٱ��r��UsZ�ګ��r���y.��n���]��1b9�AE��5��x�G79�r�zzk�uc�k��Uq����QY���X@�D��F�R�4���5���=	m$*���d� ��.OR��p!��8��fE뮴%c�q�5n[������mz^�W�����A�1�����o�/�s@Z+Q�hƓPV�j���ux��P���R1h�Kq	�J5uD	�P��5W$��&M��ƫ���1V����ר���WbъѨ�W+q�4��qŴBD��D�P42R`��6�|�6,HY7�s|ʹ�b�k� �-q,i@�t�HZ!�Z��Z��%�.��j����_鷋W�܊���Uz��^��ٯa�z�v�ͤ���X�77!r�L������û������:9��b':wBDF0H)��l_�-*`G��#��H��DA��2S1� 1c(Њ��c�����D�A���vth\�����ٌ�Ub���I!%ZFU�A�$a0�������I�;��l��;e�C��ι�Ӯ�]�`˻�Y�\#��UT2YFZ�)��cr#d��Xd����O�%!���B���UI*��@�QRJ���r�A����a�"խ,*�+���q�)�]L�a���Y�$�vx������{���ݥ����7.fyLG7����}��σm��ǙY{�V,.�r���[��x�T�$����R��m���=�X�y�3�e�fM��$�x��o7��u�I�]|���~����;E������}���?����6�;����ڄ�~��q����bIw�O�^�ޚZ'�z��������5[t���ķ��_*���A!í�'���/QԹ~��P��ʌÓ*����^(���0	�џ-����}/����iTg����6�w�>�z���|����3B�(�pA !�N��RPk��]v�Qܺ�]Gu�]wr-Ӻ7E��$Ps �D�*A� �'R�V۹v�����j��$b�H#G	FC	b���8bL����"���.�.]w5�%\L��t�U�㓝���#�M;�NX���ʽ���x��$���	q��A���S	PiU��\��[zz��f�W��;�1[r�6϶�^�Y��m+�U�^1�5��k�����$ޚ���j=wZƯe\��=���y�^���J��[��*5AF����6��������㖒��Wwh��ۛ��U�[rۛc$Tgq��(�FѢѶ�Q�|\�-��W��/��o�{�_����4r�D��QQ�S7�x_���8��N\V5��W*-Wε�V�lj��[�y�5^�u�k�����������U|��Y}7^S۶������˷*7�娌Z9ln�5F-�Qm��{���ŵ^5yv�
2G�ʒ�˛�QN�ݕ����o��6�5^�^˚�-�-^��m�G�޴!�������t�h�:܈�f%�lU|�7�[o��n��]�P�2���.RW+�^+��M�-QX�Aj-DdRB� ���&(�wW4������9ˇwA�4b�wm���E���EE��eߕ/RE. h�D`S/Y"6���<Z������^"�k�^5^M�-�r�9PA�B(ߟ���EE]7|����7B�]�d�C���)-���T£Z&ƽ�r���`�s`+�"�@�e�o�x����sW5ћ�.Wx���J���kHB8���� 		ˈ�ߒ�i��nk��r�LIbJ�9�Cv�do]�Ȍh�5rJ6����Ŷ��U�V����k^ֽ�,F�sEʮf�ʹ)�4wnE��X��v9�H՝�"�ڹ����6��U�V�Y��d�!T#���&8��J�>%�F6ǋ�wd*� �W9��F�_&�F��ۘ��ܬF���;���A
��\��6���(��s�׍x��)݋��,d�BS)����-.
�	��)��LL�KƯd@�J�(_P�� _.^���J�c��M�}]pʊ3ήR3IS7s��b	�Qb�o]��k��Q"%���EL�*Ȩ7E�m��#�
����^5��ú�h��ϓ]��H��\�^����gǹ�I� i<���t�/��e���K�fE�#� #"-��M^����U�X��&wA&j�4&"���ӛ��i)��'w�����r��Q�u�u7w=wb�Q��O*�(���S��_ �D�����b����x��N���t�]��(�JA��;�d�N\-ݺ\�6�\#�
w_�b1l[zV�C�D[@D,�r50��!%h��ھ�]��B0h���݂�,F�O�W"	@^��{�&O;t�C��we ���d���`�	Y̊�A���FE��h�'6�6�
�[�۔���yە਱r�d���망s�v��'���:��h�����	#���^wCDo�[�ڳb�A�!h(� � �R*\��m��-nb9X�Z��w0+�,���m��i�;��K�	ϥ��g\
�v)�I�ŌF�Q�h��mW<k�Z嶾m�k5o�窊-�Q�V��\�9n���wù�x�������]�X1�jwH��Kz�΢x�מy�x�	
��C	#!TS�n�#���ř�"@�	"�O���>khj�X�S��$`Iko�E��V��[�&�Tb-\�ESj���.��m���if�̨�(ѵ�w7
IMU`V��1yKZ�D�5��d�It�(��5d�(���ō�lPb��kQcE��"�Ʒ,WMc��#i!"H ~߱�<v>�(���]_�������ޗ��n&����� ������]^o�/g�nM���A���t�9�C�[gA����b{}IR�	�e��!��ohV#t%ԕ�e����1@,A!�eEG��=?���ܫ�E��y���?��~���G�x�H�_�����z��C� �����̿V��A�b��亄-�dU~<�}�cՐS��s��S^    �`Xʙ�������O�L��Y��5��dV-0����]�� ����?�UrF�ǎć���v8l)���$���&,�.�>
�3x�
��8�c�Ҕ9���_���y������¼��ߡ���d���ݷ��;ǿ	�A��W�QČ�[]*�[��3o�OJ�0���Z��/%���¬O�]�$����pVv4Dqű���{��"���0�x���Әń�6g��Y�ฤ:s	]���Qv[8�͵�V%�i8���l<���U���9Ȫ҂�&�u�kw����I��a�]l��A/}��Y�V�����`rF>�l�tWs�>�UE:p�YX�߫l�]sE�zř��^n��y���E�{3iR�{�J�R�d0�)�&�Tȶ��?���.�R8R[�;e�x�2Z��9'�2�`��ELjtmN���R�PcpЂ���7ξ��?.K?z#4	_�_�Wg�oq�:¹2+Ϸl�;jY}�<	gq�:w���QbRQH:�����O���U�Q4�t��.�Ht1ࣽ��7�
��җ�ospH�M�v�
���d�z� ���ԝM�L� �`9�(Ӹ	ϩ��i���]��6�c��뺠���G�\;�[�fL�VKޱ�֎��T+\�3�T�+9�rvHC��B��٣E�]G����c��dS���ķa��i�(=��]�<J�#ŧe$���<93���|�(��>���'sq-SW^�rg�Yq�~�q��3��t``���<t.>~R�IgcN�j�����8s�ME��T֠ɴ���L�L[���c`-��m����5Lvb&x�Lǚ�g+���n�29�?���k]�1oM;b������o_�s�����u\�7C�LRG{��Xv7cwd�����[�<wp��<]])ǧ�5�9�H�P�Ș61mL$xs������M���:U�W}�3�iXn�r�X�&�5��;��z:s��[��� �:7*m�	�W��x��?C;�Е���rDZ}��EW�ۋO���y��B��P�>���<�+v���Vu�^ⶒ�p���J֟wJ2C	tZ1[R��=}X�{��b�#&&ِ�QZdQ��sY�����������d��kM�X:��Y�T���miϼ$�t�ޓxg#:!^t �#�-1��0��C�u��1û%݇:�4G�#N�)3��?��z��ɇ����<�����r�=GR
��n7'^�)M�9Ѻǳ魩[b'��3��������`˲����*��Xw+Fs��^�<K���X��j�_0B���ON�T"VJ�'��x�}��Yr�HF�0A@�J�)s��Z���.d(-fD{����f����*��,]k�ֈ�~�[".�d�Q�L<ߧ�G;�-�.�Ա��c ���]�72���3�;s�N=�.�ѣ�I�ܹ�]��e�L�eә�AJ��x���`X0�((��5̎>/��x�|8�ݪ!*L"�r]�b�RՑ���r(��q��̨<����ᰇ��m�,����5i�[��:�[�4�^�_������S�u1F�P�޳���Q���?��;'��{�_�+����D���!����`����,��M?�d�č�p����z?�A�����I��-|�N3�A���~`�<�q(�����V }���R��(z���i�{���	H�=d�<SJUp
c��Fu�X�צ�.�Ɛ�^��*τ���#�pK�~����BL����41�*FH0/H %���'3l�8*)	�q@1�6�����\8$���^U3!�\��K0e8̓]Z�a�Y]0�s`%���>z'c�\AX���+ΔT�6:��ze���D��Y����#��g5#��@���Tn�)f�V�.b��As,f��[�1�O%�� �Y�s>՜b<�')��<!r�L���r��E��|�H��k��s�z!��1�Ѩ�4l	_B�����PS�(�$T�`B�^Q�\!�m��QA�� ��b�� ���4BG,5���NL-# �	8����Q�rH��ew��A�j�S�hM/s���o64��卭�T9����F��w5wb�4q
C�X�%�SA1d��B�l��\�Ƥ!�G�Y�`��#���J1dbi�LCܚ�s�	Ԟ| �-E�8r\��&>�\.9CBUF�P`���"4pwI��a��kF�~�a�,}Y�1cƭCAr�d��f��+ "Ě�0���q���z_6�fkc ϽD%�Xr����*E�{#Q�պ��F�qD����z`�����"$��k��"8�9��;(QU8�[��G��>��JL�3*���9i��أ4�4����٩��i�F��QJ5�o�{��P�7IH�2�#[Ed!�(�SNbq���Ѧ19��x��r���%�����p��qJ���&���,�I#" ������T�M�Nˮ�G�����'��y�#s��?������~�2ݡ?�����Rg׻������g���̙2���oSw�N���y{;؀ [S��Ώ`���V�[��ʹ�ʢ���ۥ�J�)ۄ�Vr���h5ͺ�&�e3cF2�wqs[�;�LSFɲT�D2��4l*�:�X�JţE���Q��*+`�2TE�,k�ZK��U�nW�6�H���w�����]�z���oi�|�������~�5��=��ky��;��}g��;o�����A� �r���gU��OA
���� ��36@c[����U�jվ���5kT2(Ȃ� (����
*kjѶ�V�lX�^ߦ�]��� D�&H�A�(_ �Q�E
��P�Y�G ,D��HRq�|�����[�~���z��3��:�0����e�>ۃ�����^��}�|������,{�t�`��<��A� �餁���i]��/O��ϵ����(�ݒjH}��p��(S����  �����#����~�[v�۠��dF�g9E[R�
�brT�������=������o>g�Mh'$-�Bg6;����98��/u���"���P/\�I�=A��B <�ׂ�*N٪�BEn��s�=� M���D�/e��=w> �Їdq�v�,���/�ًL�IKNw�iHpQ���6J��!�fQ-2���!���xn�o�tU����Zǅ0�4������$��-'CC�cac��[b�P#�,��ev�f.�����xd��l*Id�d��Wk�ӧ�1��6?��
<�E?4�E^��m�Mt����`�*]4�B����bt��DvV��V�3���Hѩ�:Jv�����L",q0=��a>�3�C�T��z�G�Hv�@��S�ڬ{Cu��d�X��
\��q��<����AXrb�z�e^����ڲ
j,�z2��TS�g!-��Sֽ�$[77ztY��M�am�,�*���I��#MdD�o{D��dy�P���Ƅm#��wZ���d����y�@��kp��ԏk	���|#S#H��R�i�2����y��s���zq�:Ʋt�W��w(� 0�bPx;+�h<�Cs�)1&Xb��I�8�廋�f��g� GC�[ C'zwю��O���u��}��*y�E��z���$q&���S��x"�tJ���;���M���˕#S��~V�i�'�WH0��K�j��A���^�ɂ�po�Pڱ�W�R��]�������o�A `�ԤLҐ��>K"�{���]U�_+�6Jǎ(˜[<]CT��y�-�Y������ ���
�L(8�\$e��)�$\�%�f��~�K˟Fi+�3��q��[|Xӏ�h[��9���Gy'�p�s΍����D����w��N<������AC��'`~�d�tr�\u�j�\�H�p�9�7S�뢗�k�4L*��Z+7 A<a�)ȝ�Ó�W�=���l߱K]���e�b7^�����f��<�u�N��0��m�3����N�{+6�
R�:��2uԇ,�t�u��NT��a�#u�}��:x��å�;km��IA/�ۨh��%_�[����t�S
"�G�Wx�YnI�^��!�6Usͤl��k j��
�
q��gZ�:^�h�D�Cߞ��N�l�@�x{��_���v���Le�	��
N<��7��[����|����A_1�h.{��ǄX��-���:�%��k��D(�4��5�D��媝�EI�-��s�*7�\t�=���ʹf �J��"8;tt� �������L$��G=�P�'	8�Ķ8@�r���]i�[�\wv^�\� �XJ۶{A������^��%É�pb���6c��g��C7/2��%���)	��[�eD���c�1ⷶ@y�b�U�+4�B,%*&1���_Һ�l8�S��31Ӳ�뜄� ���xCH@!�Y\z�(Cߍ/[̺�$�]#��vC^����yK����R8���λp�v\���pϊ��]������0�>���>u-�\�Կw����� ��c �h<��\_`���Xt%ɯT-�'"̂qJ�9-���p�젏o�(��x��z�Nj�kvn�w��S��n|��/�ny7@N@#M��y�=�s��˒)y�d8��!���}��ѡ������O�Z���z1?,p����|����>i��؍�� ��������((TÍ_!���M@��?���++�+���ϑ�B��c>�0rBu�8d2�c�N�!�A.P"�|�q�@No���%3[7��,�r��Q�3-�"�I:�!M8!� ��Ú:!Ή8c}m4".�m�=X�b��0X� z�$�пHH������ ٙ���Qk�`� w�j�����GV|�x��\xD�rQm�չ��*Gļ�80fŊ�[�Yq�a	$�+Έ��a�?LMƘfDe�i��mT�T�#�"�����"�;5����8�n勘2�+*���	֘!�p0��.̀�FL���mް�B����4q�,0�Y$ύ\��ϮX�P�G0g�ɷ^q1���I�r��fC���h0�QD
���^������=�ϙK(��.x �!��_Ӷ��J�|�u�X��Y��F$���qG''�`.H�T�5�1K�q�U����@�k������(AR�$U l�2�,``�",`$�\�`{��I�1�'+m����Փbb(w���R��Iy�>9��<̘�5!rRi�<�	B[)؋�GZ* !p��d!lA��Z�t���o��Q���=&j�
P��[&(A9pP ���NkA�#��	�?r��X:p&8���F�&U^�b�H�Mr�HU��F�Z�&	�0�r�rE�}8��QU�|J|�|�,��� �mSt,�C(�� ."#�m�0�H6��`����ֲUCX�H��!�Z�"�5M@���UM��?�T�  Z�B&`��"�H�ϝ��聹 ���G<X�Rc�*�kʶ�sL��MEF�MS-L����m3d�FY�c&x�-��l�XMO.����UD٬U�ڊ�clU�"�-h�U�Fԝ���)#! @�QQϊ=y>��7ŧ���|J�=O��:�%��.3�ht]�}���������έ�����l~'��3I��J��9�1y�(�ED#"�A"�` �(��CV�
� =TTV����Ȩ�|PQ*
28*�"DX�b�U �9g�����_�������W��=A}'�!�=��~����>����g��]��z����|���|/=ϲQ��_�EEoe�Z�/���"?������<�  yy&��ܔ"�����+�H�n�5Kyٜ�"���4�#�(������y�֭�[^p���x�D$�07~'��U�ό*�����׮fu�U�y��=�ڥ��L�)��{ O��|�א�X�����U�׻�`��U
�M�f���5�&��+�Y)>��z:#�E�nVך��~���h�W�ڳ,y3*�m<w���#\tY��v%d2u�'��.KǐL:�:��*}�Ę�#�ȼKw>��!���N�i�K�x|�X�z��OLܝ&�W�Uy�&�����E�,ǘ�K0��6�*�.f���I�m��]���6ƅ-so��N�����]�3�'�("��cx��\@h�Q�}�*"��!�u�ؑo��N�Wl𠽗o��5N�$V��P���<�v����|��X���T���n�-ۄ����#�����Q�M}�^1{�hS	�]�xfW  ��:�9�Eձ��a)c�GN	4Q���0iC�.�-�8�M��z͙,d��pߒ���$ů�hڗƔ�A^l�u�-p\4hL�:�ٖh��MV7�w��Mԥ�F����b(\��*w-�9MÄ>;�Q!�����8����Nڍ[t�*񺀌Q�w_��a��,M&B=�5:ո����Pu���ܻN�$�5��!j]ݟ��~�tM�V�(ڃ����[��!c�,K�Q,̓mɦլ�`��|�Q��)vdH�ӗ����.$��x>�+eCx�ץ���~R����J[㮩�DDz�9Y�7!��0���U�����,�������]};Ab�eT=]�x�ikR�H�&L�L8�4$%IB� �gc�*�����X��x]5#���g	�����!/�p�h\ȶ�}U��|���M��b;�\"b�](�$�5�f��k�9
�:|�� �������IX���4)R���n��
W�@��=6�eByt�B�� �/�I��y��KϽ�ӏ5�b�'��)	�Q��e���9n$Zc�^ojWl��(9�}n��L^R�m"~�*���˜�c)V���h:�\JNa�0���_+c�h��4�&�6p�i���!D���2ܩ� ��%4��²W-~�uRM���I�X�Gjnclӄ�d�;�A"�����̈bJ+�=��]�ǚ��ƪ|�tpW��x9�t��¨G@�k��4t�#`�t�݌�˖�l(H� ��q��-�`��D�1���Y\����}��U�B���Q��G#�n�;S�o�Z�t,���n��=_o�8���J:��5o�1�/��[ԓ���d�Jx��JlG�:��%�i�����'��{:�� [Dr��F�3 KI�^ӳ���RX�Йd��L��Ԅ�����ɑ��q����ۈ��!\h��u頺�S漧��k��[��9���FMDM�(�QA������.O�5��B���i�:����xn�K��L݆�I��G��[�o;�!�*EV AA#��x8��|uۏM��<����'��_���|���{G�� y�
O��i��6������)�<�!��*�.� �D�K!e�ɖ�J�N��)t�=DP�'&?=�S+�PO��NH���i������<Ak�?v1G1`(=����6�Ѡ]�]���p8"��\$f"�9CLUhH
2	�u�+X���s��/�6���o_G��׏���ԇ��~�A�"��׶�tH<��&��5\�(STRmЖ�  �p�)&`�J4o"��!ٌ8�j!"�j,pi�Tℸ�����l��L�ȹG�U�dTF������{�L���xA��Y	���,��LYF)t�)�ZfrD[�h�n6H�H<*�Ŧ����)@Ibth%��4
�&�KT�M	�J�N��}wz�*�0���+P���4*��P��\̝X��S��m��jF|����<�.:�a|��4�Q��T��&��	D˂�؀.D�""����%��}ǲ�H�QR�T&�`����Ѐ@�J���F+����h�X��jKB�m���R,b�X�!�Ai��L9�
 J��4�3Op�@�)�Y$/��j���Xa4�d�B�'--�WHVܨ;ƚ`�DU���y����Z��lҢ�H�f�$D�U�?i ��j�R(���1#t!�۫�%1�T+R����j��97�=� ����#�Q�E�9��V/)e����x�������«de7_������n�N�'�xHS�U����_�瘓���~ ��dЌ%[83�S�(K�&��E��?9�o��� Q�D�	Swu$`�-����hD�cV��-DmQF5F��b�WdP����C����'E�ym��w_��}���{�O컟���_��>���~'�~������<G#�v���������z�<�ƭ/T���������t;�+��D�vq=��|������3�|o����o=O�`_��
���\<�yA�?��������"V	o����L�rx�W���}��&fB��j/i�  k���=BE�?�����C��)��`���1B̷�/��_����H^M�5@yu*deP����@����N	����#"��!�n\�THa�GE���ˬ�Dun�5��rgq!D`��k�<� puPP����e�ډ�Ln�k�S���v�j�����ҡ�����ș�0K�ƕz#�YPyq���B��A@�^���́�k��v��((j-RT��|l��M�W�^s[X�;z5T�Nd�$���zpQVA��Ɯe���8�2�F�J�E�d�����7���[���<�K��i���ێ���;W����~vq�鋍_�-+v�	�I�+�[%�%HA�2<x
��F�G�����e�Mۨ7��7Ęf]����K�IC+�(����u�͕I�Zv�`T���,�$��ʕ���˕�vh��]k�>�̼��s;Ӏ�XW2{�H��9l�q��+����}��ǘB��Ĝt�6xɭM�Y?�=���e����FFKK�aZNH$�YDL��j�`�0��r�����5���I���y���a *��/�#��=��n��⺱O�v�赚��4�+2J���]��0v��,K{�.�V���\F��7j��� }�R�Fx�w��6��Wn�ap��S�S�2������6��b�5�N��b�{#�c<o��X�Q�㑏�- �1-9�udᬔ�*u'�Z��c�HC��;Z9�R�s�a�Nh��d^rO��@�!Ր�$(�_�jA�d��*u���ρ��,r�񭏘�#A��XQ].ʈ�>��!諜J��U�!��p��p �KCY
k��(�J+ݬ�fF�AJ��Q!�����-���F��k�H2���ƀ��">��!��<�:+�P#8xB���iq����>|�DGGι��#�H�;j����'��6L��]F�
���
�(	�j��s��o6
��/%��{���*6z�+���Fg���,�j�J��`�j����m��e���桌ӣ:��:��ɳyl%U�(֨����J���]��$�ꓟ2��ر���S�d�3諑��y��I���'��1	���$UX�:�Iv�D	KF�Tz7�q�����Xje��`J���L��习S�-Q$�p��x��cD>sZG<�.i�i���D��!�3�����8�i��#�s���5��`g��DgmC�ޯ@
�X�Ǻ4��1����wV�n��[�CF�!ߤ+O$��ʸe�/�g��<�Ǉ5{����W�#�h[�B�Ǌ�'y'��[s=Wtj��-�kT���u���Hu�$���u�$9�_.Fܐ�URT��%{��.�$� E�����Y�NÙ���b
>)�iY�~!���j���P�3�����C��)���d�$Y^��yZ�w�	0<5��X���.�{���i)_��v��mƧ^|�ޞr�U*��&6�G]�*'cԟh��sor8�9TU0���Q�]9�k��YK�
a�j��i�*j���b��:�S@��z��Ff&&m���;�tJ�W{�t���M�
"��7� yyZ��<�<��>��/��E C	�O����4�7�0>Z>�Q�J_<r�X���=��UCX�I�TI��������}��a���+E	HW=�`0!�P��kl�c��l�rN'���p�;�|ƣ=3Iubb�%2�m+�JiEUD�#)sR�4j?9�g|��IgD �wa�&�H�T��AfHF	ӁU������za_j�gy��������?K��IK܅�ȅ�%��V,�~�`�@;���9B���8dUL���ԺC�!�':�zN"�-�Tc���T�H���CS���
,��/;I2�c��A�T����R�]T��U���,��(�i��-�~�|�&6��2o�s�Ɵ�K���<�=��;�/��O�~��n���a�~���߼+ӎѪN�f�|�ߑI�֌r�C�*�R$�x�hA��D�H'�b�XA�0F�"=E f� ٦lWJ0�f4�$*��[� ��@y�J�h�q3��!�?'��o^�m���5e��m���{E��S;g�o8��0���nM0J�����H�'RxA5@��H��=5��H�//ʳ�_�~��|�C�Z�/q�����}0���������$枡�@P�&:d*�>TʑHJ �N+K�.�.�	~N<�m
Ĕ��$@�P��	hN��Y�&����4�U*���@�@¢Jl��{J(H먥c��xPU���,D-V��1]>?K������k�Ӷ򿯬�p�R��6s�� 8uו��WmWR�H5�F��V1��<4��{�+��$�Tj��ҍQ)�4dƢQ�R��5�v֡�b�j ��m �@��I )��_����+�x_=���7��ݟ��ݯ�v]O���/S��N���{�|vg���w��~��w$M��m�G[�1n�D����Y������4bj���IP:�t�N*�g*��J
���2+��F�ev��D�ްx
��ɚ����]XhL��J�Z0s��$�[u�
̺��Qfŋ�4�a.[L(��q.ú�*�]���3��꾥�u�˰d���bR�6�Lٚ����T!x������WU��8�*/pH7�]���,{��WR�&n��,_ǡ����	�1��>�.����=yU�q�Ӵ��D�i;�
�VlY��Ȏ��;ӽ+&�$�{y��2���obH��2�r.tV76'S����Ɏ�N$��"������;�Ak����.M�A5>ﵝ��'ٞ�e�f�:���"����mrD�c:�!d��h�R
.��Q��|�V$�֧�v��u�ysշ��87@���cf�[�2.�]���9���ۡ�0�+�"8]�F���uk���bfa���B�n�nٻ�����4���9�j�[V��V ��9?�r]/�c��+��ngK�x�wN���_t?��>��t�G}���ꗹ��If���������>��`�?=f�3�־��5�u3������17ƅc�O�xW�<��ٻ���p��-,/4l��+T�K0)+��sVC��̀�>���e�҃.������LJ�M����V5�~��{lҧ�\�q��A����t��˟x�1��.q���<W9��op�|;�Exs�dѴn)�ZA��!��38!?pX���Hͪ�>t!�
�ʏ2��tn��)�C����N���#�%���b�0u*��,T�;n݋�dy(6�gOڇɀ���P�,ܨ�	��1n�A�JS�X��L#�o�]�ڲ�w�1��������S�w�1j;nn��pe��T�&C��۶�Hm�����N���M�	]�|1J���gq�␏��ǌ2���X�[�5�/���to�M�?wC���Q�8��dh� } �)QA*'�Ȩ�T�>r��!"�saf[��1��Y�'������j��<%l�N@�Ȳ��,��Kl�VZ5u�,D��}��#�?l�gHF��9�r	����@0�|B�!e�]�Z;�Ip�UX�d��]��Z������L�߽+x�D���[ON9 ����N�'ߗn�B�*N�K;����4z8��k�lϛ�kG��]�|>�����Ʈ�%����=�f1o�Fb��XP�Q_>=����6u�!��x>c�ܸ#0b*j���AO�mG:����?���ӑDG�Jb�C��Qi
�m�� �g^�n2��*�8�Ν2�O
J���e�9t��*qߜ�Ѱ��ˊ���c�η	�7�u-H�б�v�@at3	��`�ֻ�"���W����[�+�{�º!�N$p%g���)+u�; �,����=�;���:n�eؽ&o����r��p��4�#g2���ߖ&�˜g`�cC�w�n}�+��]�s����K���%�&��!f�]��:��nkĜٛ�W'ٻ-&\g���� �93�XZ�',���d�t`��i�<s�����$�7>��4ۗ�[�'1v��i���u�=w���u��6�%n�h�"�������ꥰ�ݫ
�˹)my�>����ܰ�*{R���`�����i,����0LB7Z��y�p%����r����C�a�cl9�$���#ߖ=�5B�!$ʧ�;�2�p��3���*O�y"#��	Ĩ�7Q�:���ۂ2xլ""��I_���F����PiٯE?�z�qV�r.�R���U䌤��|J�rjK�W�ψ�f��rӺ�6���I�֑	w�3qC�z�8��.FQ�v��;!pf{$���r꼩�̉ ��/�Gɞ3Gygj�8�a rQ�ےWT�2������t^�ٷ�bp%E,�W�4zٝ����:4��E���:d�`�dDzc	�&����'����b�w�$pC�l0�MG��|o|f���L/��.��F���I�'pP�zp+lF��g3�w�����"���{�����/tcwL7�֬g�3r8 s���u$�To�"� �9Ś,bm-ܹq*�sF�;-�9G��V&D�v�D���y�jm9U�OL�od����g�l�V�t�x��+��O���[/!ٌ'�'g�!�z��J�3���B?�x�p�6�8� �>�a��,�~�,�^�}	P�C��^`<����?_��уH?}�����B��A��y� C���~��AS�@�C�=�Z�dAF+��Ǌ$6���I0%YeVK���$�XuU�].P�d�xK$�*y��ހɦ��.#D/�̎� e��1"���z4�ev4�,S	��t��u��7総�_/x�F!n�t���r)L������������Z�:���e�oo���yۻq�O�����͗����aP��ɱ!,��#
H�7�x�EHc�M#WP�n6 Q��^Yc5�[x7�"S��J{��1
��9!l+9�AG���Lh!0dJ�L�U�yL'ax��E��R"H�x�Sz��$ꁽ	(�:#���	��6���/0��A����0��6]����r���ie��㟞z}�=�^^_��}=�v�J�*���۷I��m��m��A��X]y_>��6��[������$�QA�eD��� 2ǘ�W��}�fl�$
e0����[���ɽWV�ͩ9B)o�ۦU�<tG��`�!KD�S>�0��Ɩ��@��0@%&Y��X�#dIDI�C�F�j��r=��x��j��^�ۋ������w��|��~�8BO3���<��(�00�í8!���.�T.��۰���N����^;�/���~��_�7��]���p$y���"� �<ތ�H�$ H�V,Y|˰گ��i-F�n�W��!b�dI@$|t������bw_��dUG��y�wq�>?��|�������z~G��[��y�?g3�}w��|���?Q��<����G��%��7�����9�ܸ�]��L�/+�4P�D-M�ɍ:''�!�����Vc����N���Mȫ٬AEFȅ���VH�
� �0,"�;s��%�Ó���a[1)������9GU��YQ�s'1��Qs�(���ȩ���ٵ���nr�R���؛i�t�{��+vMJ+3��z"�����<���܍�!���:b=b3ΧV豑^㍺�qJx휜�ݣ;#�eFI+(4%���u��:�LE�D�ލ���S;��(�';ޡ��=>��G�JE
�E����"�)���"���e]j[C�a�lo;1�ZZ�jቓF4z�}�f<�L�fb�W��f����q{:��$u��Eo�3{�fá��k��9/�_�C���&�B�OtB��k^��{�<y8��ZS���D{��E=����oAc�g�֘�7�v�A��7����QV��g3;�!�q1�|����Y����f�Q6T�ϱ9����f�T�O+�9֮OlEr��]�h�R�M�&��¡��alb{��w*{j�f�gx����9��ˬ��@��_N]w\�经=��)1xyëǕV��8e
��$͑#ג鬿E:��}zQ��LM"��{����5wY�vd��*���wf��
�n�5����U����;�0`�ةs�0Q�'&{�p�=(��=Sp�q�5pEi��Ʋ��7)N.#"&fwS4&.�wSeK@*�t�� ��o�/��?��ܑӗ����=�=��_RyF[�������T�}�s�|/�?ڍ�#��щ?u�E'�#�o�
X��
��\S䦰2������ly���f(��LtPS_� Y|�	��W��'p �`�}���@�|�J1�x�������7^�Y�m���F���f���9L�A�ẽs"��*���&���{���α8�@�ɞ��R*�ײ��2���.��]*#���I��],��P��D�s	t
�ߧHz̶3�h���,
uO998"{Y7^���4
��#�Q&i:apۏ��i��>s>m�"�)EFVa1��#9и_q�#�;�yuk�5J��'r��&%R�fz$JS�Vd�[ *�n�H����x��������x��#KR�����ocR��x\�=�I��^Ft΄���+Q�F�w��Iu��� �l���;�g�%�i�	�Z��r����,<r��l� 7t��ТDz\�%}��i��C�6���fv��tZ[LM�k4�V���qk����.�$�Lq���e:w;f�Hy�^�G�eT	
��~�=IPCw%QSm�H��m��5U���l�W��i�G�lh�a>�f6���$��QkF �^a�V�E8��k7�a
1�r��Ю	ْ!!�F��u�j�v�~��k��o�L�W���"�K��-�*W�3��f�N6���䰯c��[9�������=�{M�ӵ�n�4���{�q_~��夓�����!GN;u8��}Q!�]v�h���ش^�8��X��lpٞ����o�Jg��U��96����:�:{F�i�4�ӂq�&�B��Ѡķ(�v����!�[q�WqA�S�u������(�H��ǀ���͔�����K~e���p
ZEA?�rSu��z�b��Զ��^��T<e�x#�0������USQ���75�-(@�6�`bwc�oS�$M�;ld��}�6����1�)�#[-х�qC���)�hz�=9>��w"q%Rw7vL��kq>b�=�ǧd��uY8�o0�+c�N&�Ŋ�ql�n
��5��s�AϺ]�p��I-tNݻ�-z�՗���;�ov�3P�ѕ�=���8|tPL��/�N$�Jq��)C���#�`K�n�3��˵[*Si���*��M;*�܋�N�ܘm���WiZ=B}Iw� ض�y�<i�u���ֻ�GP$C-*=�;���M7�]g��)��7���Xl�r�.����4���c����rsd���?��2q��'�M �©*��	,��S4�Y-�5+FF�M�S��d�Q��j�5�a:��0��4[��E>z����)
�	�C�i��x�ȷ��I��t/�C,�%��,D�^�2t�xο(P��в`��
�&Y����[u���r��It�,��j��"��T'�x��¸x�`RI�ǈ�pdoUm�>�$���� �2]8+fܬ��
9�>-߬�#�G�JG\:u���[�4^?5w��e��:$9A���'��v3aG'9E�v�ߨ��K���]��ъЭ
s�
��@��N�#�!�
�썛p��]Ew�	Qs\��'���S�k7�����|��W��[K�ܛ��۸	U��w�y]禿��[�y>��zmr>��x��K&}���n���kZ�B�;�=4۟��C����/����o[nF���S����v�?{�_���_�ޟ�������_�?:uH+GZ϶<˷e�gө�=�J����;���<�{�����+�Ęhq���i�$�!��}v��s��ސY�	��5��*���1���X�S��z��Җ���b��ӬN�^'��یQ�}�����/����O=�q��/����1����Bث������ƹ?���
���-q��1�n�~;v��~}=����\�Ǐe��m�u�xy|�,�����r����ǯ~>g�%֝i�u�eox�}��έOo����|t�]�/�����>ca�o�Q���zu�=_�L�7��[������P���3���ִ���M�^����[߯	?j	��vy����>��3�_���t��>x��oc8k�ོzV��M-~���{2���!�r~1	�%�M��}>{Z�M���C�u���'��n���}��ti����<�K'�>mJt~�a��i4���
��I5��)˜��Z �V���i5�Ō�T��؊B,�H2+ I����m��z��o��7�C��]���_��{/���O�����t^'O��6��K��_ߋ���N.�mCm�y���x�کa 鮼���W}�8��@���e�2G���?�I����2��d!�Q���Dʔ���B�$E�&� �f��h�Fb��.��p뮞��s����ͭ ,�,
�X������>2��:ns��(_��=�D�������|)�ɢ O����{��{�~��U��)��}����#�O�9�|�R�%��{�ө��� �|�|O����<� �<��:�n����IR�����Q�C���tӧ�����N���wyy���[e�|�>����c����8h�[�0\@��&�i����T3ۛ��dmu�g��ҠN@~�(g��<����yy������������Jw!Q[Qt���2�d�+��*T��\!�W�V��r��a�~wa�0��>DC+��5O�M�
�����Q��e��B�� �.s#N�GdTu�������i�\혠Qn�*�f�ȟi��^�7À�:Ӹ4�ĘI�p`�s�ʽ�R����񰴩̈�K-�]w'=B�r���j��;���x���%ȇ�	���f�n��|�8$V��Ù�<�cW�h��ef�gp�r�]�Tq�!@Aw�D5Fw<B��E���r�Y�a2��f*A�V��}W�3���1�ׄ�������Snwy��G^\��-��t��+�Z+sl���8c��La�8
��C�=j	Dx66��?o(�X����cq�q��H�{ �L+�i�1��(�R�=����9+��:���'.[���P0�v�MlF�+�ġ�ۄ2�j|	j������P)ۡb[4�y�v�P�D?$��d��F�/Zh����%v�V��,\H�P���L��G������󓙧(μ��|ꭒ�C��כ1o�`����2`�,�>z�5#�D�A\c3Q��լ��!���Se�;�e�xq$ޜ�%W�pl!ߔ r��� صX���M���H�s�v�Piߓ���L~;�٣y�#?Mq]�59���p�A��o<H�\��%�8�K$\K�V��6��F��S܍�̵��SHh�1�8_��Y܅�w1��<p�l���%ptޑF�6��M�f���/L	����G$4�s��*u�W��K��%�3���#�<v�d�	4�@�>��yS6$w�1#�e���wmA�jg�~`�,���:	3�I@2��X�����0�Ѣp��옭Zx,���M:B6UTը�:�c(Z�ZԲ�(�w��S�crQ������2�w����
��Sk� oU��@�G@)O͙�Z���]y�y�����1��~U�'6jD�m�5�d�ӏ�V,q�C��,�	�1����WϢZ6��&菂�8�+��q���gRU�Z)�\�Q��&���sK����M,r\8r����)KF�[#��8��=$�-P�$�s ��|H�U�.M��P>��Ô�2��Ye�CBלR	��ZUZ���P+;��h�e��;�s�8���+[I~JT�!B҈m45)\�k��<���uRVdw�r�:"�ӼEg�+E��zZ�6�ٳ\q�X	q�K���ׅ�6�mE7�W^?*Bq�Vs�0���4\�ţ,2�O���p�eU�8)�P4�6-�S9�@]xO�쭵T�ߝ	-��ӛ�mN��I<��v���s�i�/K��QMf�~am�d�6�L���%�z�b��;���3�_1V���+2Y)aծL�u{��r��hi6�F��t�f����;�j�j�w�H� D�N��Le��E��x��NV<~8�N�7*����������:K��AD����j���W�q��ĥ�)����=���}����!�H���]����z72�Ӧ�u󖿿T��>/z��o���n1I[�jx�zm�9.���Wx ������ �qYzz��Q���z6w���OQ���5��<��ܫ��5��4���q��(��2ڑ>=2�i�v����K�~<&��t�xѹ������m����H�=�e�ԇh�:q�t����A����[����tZ�8�Q�=[l�xno�:o�D�m�R����J�)m��x�=ߗ�i��~���=%�o��}o��[.�t����Ǐ]4��'ĸ�o���{S��i�Ǒ��8��`�4G���+�K��\פ�g�<��}{��ﾷ��z��<K�|OƏ��~ s�/=x���!���Z����񷬽3�|���?'HϽt펯�7�ֶ���7��s��}Wpq�)s(���zH.����?��'� � FC��x�6(L$�H�$�HEF$��~,ݣ��y�5��k7������\�G������z�������~�S���y��>˔��ͷ�w�+G��&���2���'m������L�W�#�"�69��y��yw��&!�[���+]Wތ�o2��h��ک�[���;��l�]J��E�u�ctL��m^uE�,ӎ��U�,�>�{3�|��U`�zI�]UWϝ13v�9�مq�W,��	�̉��6"�MGfL�LV�<�.<�]�)*e�u�����i�۪R���)^K�4�U�éVLNV�R�%����zf���A��m��P�%]�
��	�(Revu�8�"����Ō��#���+}j,�%���u�y]��l鮊�׏V,Cg��]7.��<���{gkƵ�ꍮt���MN���4�(�4%ND�k{�����]]5'mܜ#R�Ƀ]Z���.p�Vۓ�\��Gb5��_D��,���P�`1t���3>ڧ�V3 т�DtLs["UP�X��r�&�"�j��n�#U��Q��U}�*�动h�1.�]b��E)��a�_w��i��D͡-:��g������6s��e\E��=?�Y�m�9���s��N!ͨ޾�Ȋ��),�W��_-P�ӳ����m�����Tf���sq,B���f��p�IS��D�P:��$����I���B�ӯxnf�4j'زn�WSS�z�����Y�t�:uù{��o�-�;���/</2�#��kr)��6ܾj)+:�Es�a�Վ���q�1eu�IL�pc�C��-n<�y�ruu^�����Xܣkb.:���:H�[��H�Y��Q����ύ\=v禚y�ӱu�GaZ�R=�&n�=�fAћם�b��Sq�jhvU�5|+&�&�E��ӌ>{�s}Q&�����'D=V{Q|���.}���;B/��MZș�O��<vgNȇs�"����Q�Nn�+l��ww�x���m�&�	���q^s��x�������3){+�H���OgDY���2�VNMT滚Y�y��w�����%��O<��fȪ�K{�>Et�Q}��¤wT�<���^����ޣp�,��ɷ�����=Xcqu:���V�V���E`m��z6���1��U�yTmwM��}ܖė�q�{�k��Z��Q��kiR�'��&�x�r�M\\o_];��s)lU8�	7�o�LFۋ�]ƫdJ���V��d�L;�ӈ�oS���V��-�:��Rʘ�r�:�tSPA�]�٪�|�ڤ��.�:�l��_������I:�]�v��>���S���ˎ�)��^�`"*��E���!E��4I�$�"��f2/�N���⛠���]�4l�^C=UC�je�0�{x��;�*��s�+z*Q�#�K;�q�r�d-̬�}ވ��zSױ#���r�S�27��n�oxN\�����'EQQ�竞tYٻ���q�ʮ
o�tB��\����1�M�O�'pD�ӛ���F��l����QLH����;��f�DY��<Dօ��7�Cy΍��J��;)Z��1֣J�x�쳓�K�ީ��d[�61�沜�V�WM�B�g�jfz3+9R�(�]�d<��:h���Bȝ��lfv�&������lÓ�os���"��O���k{#_&`AWwj�\�ި�;V;�a�4����)fj��sG.D�F&3�칓P���1�Y�}�D<����We�L㹲��/�\M��s#���'��4����rg%M�����q�M�*���w�MVd�K!�/���z��_Nԓ#��ypV�d���7ò��.���3#�;͹�B�����]�2�s�K���3*M�Ɲ�����JE
kv��l0��,uLf|ú��N�U�֨�-��7'�t�ޅtv�K��(��'�KF\���Df��]V�*��	˼8��Ե���Oq��.o"�5�zs�Эԅ֨Bf�R[�}G7th]73�*�IP]Ѧ�.T���S[�N:��c�+��lnt]ج�qDT��;L]N�]w����o�75�^|'tp�a`ىɂmWn��Y��m��-��V�76p]�.���v|���=�&��ji+�>�q�F�����c�f҉�L�m9QuJc/v2�T�̼�G�p�^L@��GY���tkQkk�����ܑ�i]8���q}qA汛dF���p[�t;�c��䛮U�ê�Uk��\nt�J�./���!3�#�!Fѡ��Z����\�ʮ��G���fu��yf,i+շ=�Â�2���.b/��W�U
Y|`b�=B-\
��l�ؖUR8��F�iN�6�4���v2h�v�Ҩ9���۪��m���@:�C�KU�6�dX�X-�񉭓��o�u��[ǌF��	!څ�惕�D�E-���ь�wa�EoVf��z3i��΂�B:j���e��"�.�ҍU]Ӯ�b<�0m-n LQ�ɇ`�h/�N��ݷ�ۇc��Η��ihsM������l����5sd�:����uwt�v.�R9�*F�L��S��KV��jkd��Gt��foL+�f��إ��Wtewm��Z���&��۞ɛǍ�ڨ�ތ.���w�gq�9�	�ȶ�R�*��iq엑�z�#u�d�L�'�S��Q�Sw`�6E�9ȚU�U�0xt�=����&N�c��]�3<��;�p)G��;S3\�&�L�Ը|
:�Fi˗VLvH�1���G;2&�� �m���<�UǗ�K`ˋ3�t�5�P����D��yф�W�{�pJ����
��v���tH.�8Ԧ�ī{5�E@�I��ێ���ʅd\��69K5U]	V�����0�)��qAv�q@�d#r��f�-r���JY�Э��ܣ�37l���N�F�_�!>9k_q��כ�Y�b�yX�c��B�z3��Kx���z��qћ�76��U�R8����5]&���͎xC�k6;:�qC�Hr
��݌�ٍ��{�W�«��8���ƣV�Bh���1���k:���3U*�Oj���}mÅΧ'5���=�i��`5�k���b�è���ݷ���t�`�F#v��L`��-�OMVд��ב���{ѕ�=�L
��3Y�^�k�[�ъ�1�1Asp"�+��ləsNA]c��T{�m��'TlOt��p��]P�.����Y��<U曍�Uvr�",�Y����mnF���NH��FnK���W�ܘ��g.b�v�%�B�7O$��s�A6�c��E�xc{�L�q;6�ua��tvSJ;$�s�ywfL�\>ɘ��M�+�;e>ɷ�˲0�3�4u��F�nUfD\�s��WQu���\�jo:KbDwv�C�z�ќ���tV��Nh�bqL�R%Jrj�{A��A��ؘ�1�Jtj�sWu��vMf�������wO=����Ug"ׯ&6'�r*��#�����٩�%v^5���6c+h�"Ⓝ5�bTtM�km�F�&,+����ް�Օ��%ۛ��o"�)�)���U��ϔl�zh^\L��P�5�w˜�s� ޹�PJ�j�\��=�c{�/-q��w�+�%�iF����uU�λ̥�,�OiΑW5���;��zt.�ƶ;]��\9w& �;�īf�/7��V�ۛ����lZsV�U�<�o��x.=�#��}�Ug�{[4;&#��^��2"E^C�3���W�G�ѓ��xt1Mɜ��]sن��M�Î�s��S��g	Q!�X΂��Sh�]j���Y�:ÓQ8��͙��f���Qb�4���Ҍ�߇v���'-u�"qa��UU=�]�-56�>Otb[�:�Q�;w����&���TSU6*ۻ7�Tz�v�(s��x�'zw"�TN�s��ي���}�ֱ6:��[p��.M�'���oq��w^n� ��It�-(���;�t�]�f�gQSv(��#v���v>!2ʭ�ᆪ+v�yΝvʰ��V��k�]���S���
2P��)JU�*���6w�]�7y��a�{nA�]�d*0��/�Wm����}�DÝEV/.��w9�͒��dܻ���Q]�ߛn�m�n^e��e�L��٘�Q�չ9ە�D���k�����$[1@ȫ�ז6�0f�5�Щy�=C{0�����[�pk=���l5��<��=y�BńzƉ	�MNN�k�˷y	���t&a�
s.2g/�������޼�4��[���WJ(�
츅Y��G���2���mj��iȫ�G9Nn�^�Y��fI��"�Ԙ3���NТDf{�A�w�#����_E�߻=K�h�4�]�Q�n�;��"�{�w.�OD�i��hW\��=2v��9�q2�c:� �6;(�p"v�h�QF=�chV�&�{1\���{WbD�e��:Q_d� �;m�:$�n����5H�،7*4Ԩ	�����ə"j�Z�4��;[UX1H��{5wN��j�m�C�i�d��^��yJc�ٗ����xA�KN|�[F�bq�IѰq�*��M�A��6����\FK�8﹑����ۏ3���ǁ�IH�����3Uu.�F�n���ڸ��tb%f1�C��N����83��(�T�j�������25�`�s��z���ܙ�n8�n}G}TU.���:�9����僕���p�e�FM{���9�;U��Ev���ݓ�\k)��3]P��\q��Ɏ;�c3�DJ1,gq��tb���5ySԲ�3���ynݠ��Do,w��I!�;5�Xt��r���ص����k�v�m�ջm��yd�dX�ʾ/iI�;ffjb��7g�}�l�8t���a�U�����СJ��W;��mE�f/0,�w��w�wgEdҘ�Z��ǩ���ǌ���M8N���Q��G%2�I���ا>d��GokER�6K�����׹S7�GoE�١]J^�օlܶ�Ȉ5�W䭪q�GbY�^téX�dS�[5��QM�˗,�
Z��Td�¼O���'��im��{8��+}�'E��/EmC�oN,h^U^:�7+�ۛ��<�QYfs��-p�3����ם�V��	4�B�4�Zuu����|����ƨTS��c�P�=���Ta�\����T)��)��gF��[�D�_Mw�nf��|�[v�NvUwu�ɮ}�4�K��ɲ�T]�D�Ҫ|���=���Cw�L����f��AZ�1�M�Y�����=�#��%��}W�*�&p�P�����ЖS�^�X��Z�g)�Dz(�N?\E�l�.��#Ab�c%9�k.t���أ.�#��%��!'�}r��u�����$�U2��t�T���]�^��6�f!����s_[}iċL��-f�d����ES̎�ݨ4�٦7���ʺ7��q�6z��i�Mh�����=��c��������|��\�"�NQТF+r*Sa��դН6ۼ���*�v;�9T��yos&�z�
;���3ul�S
)^�V@�[q��_)�v�B�m^���;��a��5�P=É�#%P�ț��S-92�u4�������XLWg�sN�q�ojkU)�5r��"%u��S��N�N��r��6���hd��w�:�]r���8�D�F����@Θ�b<�3���t*�q��n�|�U8�OD�ޑ���曘1ʍ`� �Q+/7hM=����]*-��U�
��mp�9*wn kMD]<���d^��f�f/�N3W=
N�:�SN��wA���ݕ��v��91�F�,G_0�i�u*��]��7n­�9s������[F%9V���Y9�_L����!�s	���,��}][WӤ.�]*��]��Bb����ލ��˃��Ȯ<v�!��X��dGUۂ�ˬ��IJ�wڔ-�t�f���r�.]n����jFOR����,���ѐ�gk�Ng��]�Z�P^\[�&��Qi�U�p� KR�B�ښ7�k^(܇���Im���;Y"��Ϙ������Y5qy�=�]�4�5�VH�Gy�S�ՆU�@�O8VFvtf5Qb���V`ػ�}�!t#~�[��bG�5`���h�^�w�����g��n��3�,Fճ��UT�,Z �mu��ݞΛ��X�Atv sEE�Mˠ��S���"*|��mC�vA�Bj72iOx��d�^
�t����7����&*�>ؽ	ͪ����$Q�X6���ީ�5���[�\N�M��f4��Jb�e�پ76mAգL���3 ،�8����B���[U�'̳Z��Yd#���f�=�Y��;:���t�U8�Pת��⽨ޛ��qݪ��9�����5Q�B�O�[qP�(.�<����:ЮK�۰gR|��q8�W��5:6B�6�By9m)3�F��J��U�&�n���ؚۉ��Yjb�ԉ�0��C�ݙ+�U����	-���Ń�us3s��<�|���,��t;1a�H��\��s	Ȅ�7; [黨Z�q�:���:⥉���i�Bb�Ήw��L�a"/4�eu�!�4�Ӎ�Wk%�]��ʾ��l�e*�XQ���L�9������&Z�Y�3�c�Y�@A%�J���ز�nv3�Ud���Sb���#jT�t�p���z���	�Q[ف��6.o2\�G�oa��zMT�b��qJ�\^>��2�f�t��v��4�X���&3`�����ËDe����ĳ�{�u���έ�4x�X�����jl��S\��gEzs7)���
˔��QꞨ�[=�FT15�ơ�&9�|!C�U{�E�櫺:�H��{�;�qC����	��E�.;���u��!)2��[�9G)�-�Qv�e����ip��Nudk��&o/�P,��cbLmtTv\j2�������v����"�+R��E��ǓU<��ՙ�:͗�T�Tu,�ˡ#��R��j�����s��fj�ekRѼ*���ݶk+zv#h����7v��^v�5f�T*�.��^��HtoD���j�:�L��TuYfM���ݪj�h��TkQ�dm��{���{��u�;��u\�%V�%N�fW�{Q5�/����7.s6o;�r�VI�@��W��&r�'���՗�C�p��݉FaF����jv.&,�0*�u����j��U�֠n�t�܈$�����i��ka�״F9��r�Q���p�6A
���ƱoE���{%i�a��ʳZ�F�Ԩ�{��ӯpku��+*uW�R�܋�)b��)�&���v级�M�] �����Z4nVJ�����U�9Qy�g3P���1Kv���z󎊭��/���o�AY��f򪮒�Y���=�]Wu�Ѫ�y7��Wly��P��1=Є8u��W�U���Q]�y�Z"�O<=.���6�A�kb�|^�/SO��2.n��^�ԞZ��=R�p�Α=>%M�o=��0�\��m��m	Rf���ܴ���ݽ�!J���o�5uh��}g�.��dc�^q�˚bbL�tۭ�˅F�ko�]a�/t##�U�re�E�����7�E�:v(�k�ڨ��NS��r3^��MlĠ�"���Hr�ww��Tbb6�z������WwJ�.�̒d�aop>�+-@��jҫ��x����m��/
㽜���v����rF��g�P�d>טTlveoV;�b�KŰk0ӧ�3l=W��#�vRU�W>��9s1qws�(4�6ѭ���t���0QLK;���ō��8E�65�+)�ꈍ�;k��m�E'(_������*���� �TTX��`���tX�d�V�x�یS%,Y����y�
��� ʔ1�Vj�.��̫�hMQ��Q;�_���iWVOU^[kM��﮷1l�۬)��<��NlB���xV�|4wu	t�lX��6�;���c�e6rnd�c�(S�ņ"�/T�t���MC�\NfMc�+��t@�|�Y9�a��,aR�`�De���8�u,�Y�ձsld=�cQ�]9���*͇B���vY��Zܼ�B���b��'��'*��Jnx��5w&��x�:-7���|f��n��5�ϝSvᕑU�yf�c���.�zy��/0O�����������c�b�.x����Շb�;O<n]���Z{0�fռq�}6amf��p����$[�{û�`<'DZ�:�s�V�Ő���%������D\����r�;t�P'i�.\H�SעL�궮��Ds��+�X;�2�`�jD��v7	����
�vɧQ.��PO��R��L����^�t^��u�kk�X�h�pp��SGfn"8ӂ�m�8��&��^f���j%�������T�9�\Mt�<�)Ѿy�L��u☄��K��s��)-3F����&K�uY��<B�Hx%N��*���'�QγUt����gب�j���o��Jp�9���!=ԕhو�iܡ��%o]U�٦'6cv�!s^d{Wc��qXj�.��"d��\�U�	\@����w�
-c�47���f��m��s.8��!mr�ξ��5
�{	E��t�՚0L�ȷuV �G��jTnڀ�ӈ]zu@��Z�s�V%B���s7-�ܚ�T4��+Mp����YqW9S�v��T�ZP�c��D���٘��a�m���Fz�bɵ��Λ���z��t[H�뚊�X)��z]
�t;ke���꾩�2'�WlB}f� �ړS�]=��lr�荨\b�{��L��Tr���	��j�r&����g�q����Dc�}ٜ�<)a.�-(�kay���]Y��;99mV�qy��rnH�h�m>������_
�ʉ��`��9�c+��k'ݽ�����ba�v=�M�U��]b�1	��,L�UH�,e8�~(^aj(h�ں����sf�"-Q�J"K����:�cS���;r��"�& ��껕}�t�/5�k(�FP�s���)����p���|k8�n;]:��t�.�H�5S1�g48ڨ���{�I��ȧ��Jo*�G:��Yn0�q9j<6��vL;�U�t�`��y�xv.�-ĭ'�Y���Y�I�ݐQ��7�3�uc�.��Rzpeݭ����v��s�oc9�δ6�S�R!Ld�̰�r
���2s��+�f��+*�oF�N�t)��}cd+WX�I�Y�#�e�f&��ܫ�wR���n���.�Ҕ������Ħ][�z��_�
�
�̹������5���QY�����$�`�w���*E_,��^.�m�}��E:Sәx�Fl[Ǣ+�8�|���c��Yh���T<�r�B�4�9�鍍�v�eI{�#�͚�՞�	W��f�j����;'7,�1HYr�v�˝�b�����\�9Y��teOL�5]�#u�I槗v��������]2����OWZO�pnY�ڛ��݇��b���Ԋ��5��VD���Lɚ���r28V�nVf���9&nT�����hÚjg��t��es����O� +zA>x|>���G�Үj�I��kl�)�֙Ŧ�RJͫf�Ե`ikb�lmkp�ۤ3-�r��;��[���m�ծmk��r�5t5�N�+,s#�r��dL�12b��:�9r1��t�ѱD]whD��U˹��ۻ�U�wV�si8�(�Q�E)�U��j�V&4gu��r�ċ2K].���pguu��;��۝���;���Cs�����ֹ������,h�u�$�ch�U�W5r�,TX�r��L����w]sr��.nRRssnp�ms�nsm�Q�s�.�6-�t&�Z1��Jwls],W6(�9IG.\�n]��J滝���*Kn]��MPW(�s�]��]�sj��nQ�snQ����r"�ۚ*6��܍���I�nV(���gtW*�n�5���+r�t�������"�F�gtmp�U$��+F��r��.�k�ȍ�!�V�ۜ��An���Ü6��ѣ����Q�QW��7���tרZ�pW��D�����;j�9��<�K���w�g��{~~���|wI�q]/�����~t��Z�C��kܸ���Co�9�¾�ލ�{��3�4�y�2�*�=�9��W�1����~O7d����
�?���G��6l�>Q���IO�<v���P�Ge���SK�J�!�.Ag#�&��-c֬��?�ߜ����M��,Xy������8;k�/�����K����ݱe�`�� '�v�4�cc�
�a
2���Yq�w�]�������2�W��E�S�VD�Ͳ8�I�����I7�B;���b�(�_�/-�������*l-������2"�>�F��X3�p��D�>�L(H�zm�O̵��ɛ-���+�~mj	"�"�¨�5Mh��4��M�9^'y�Lv!�ᶾB�A:����1�jt�F�d"��*��t	P��
7�	�E�O0�z-�i����¢zHp >���|�A��v�p\-�vZ����l�򽍓��ۄt+ٜ\XN��ݻf�TS)���]]�aa�U3���9eQ�5�s�ڈ�R�ȚDj�-s�r�w/sn�q8%5��3���>{0	�n��R[�⌝ɴV���Bo��<x���ʗ.�\[�3ec��h�S����4rk�!cR>:%jw�q<�q�s��FP�R��#�׷ �m�[�h�q��.�������Q�	���S�#B��J�^�\�+�L5�M�yD�l!e8��fF['D�D��۝]���0�l\/��*��v���}2�A�u�*�b�S�����-��ֶX�@	T�m
��`Q��4�CvuԈ��C��l~�䦚QV��>�՚� �W�j@r�c�۝(_��� �u!X�#PN�548kD�8��g�2>�>ȅΫ*H`YM'^=7�"�\�]lyV��
�pA�\�+�Z[��+#�i
Ȅ!��˰��%�׹1�]Y;*u,���8_��#�7�۱N��N�1�!t����m8u7�]e=C��qpN`I��De���D@��n��)9�0U�Ռ��1�L�2��Gl�ZI�p����{���׊�7C򧵺��bcw�t���/t]��y�9'o'�������lz�l��4J��!�y{T�C1L�kmH��LU�r~Spa��J@"[�Y!,7p7�)�E\�	$Wsm��L�g6����]2	��=�j9�y��T:�[�������b�:�k(� �*�,��#0k�����Vq�S�m�MJ�n܇��sھ])掂k�Gi��o��!t>�2jǢ�S��y��@�=��Ʊ�ym7S��H[>��wa6?�*_~�DTE�z����U�;)�a["�m�Gpκ���+���a�D�*�m�3| �G�&ؘ�Ü!�AW>�B���Qt(��ǽ��T�w�桝�)�C�N4.�]�Ы1�:��a��#:�x<�ύzʱ*��3Y�̢�A���J�i9נ��l�.�4�6�����Y�Q�-|xT�Pܸ�Zf:>Yg<m�oWxp���%[q����@P�T���;x}	R�Ƥ�I��p�}��h���q�H囙2���Hbb[����#�� ��ŭ���|�ͫ���l
�a)s
!�2D���lcL+�n=݄+�H�o6d�|�VfCqw{�AL�_��ã���_0  �~v� ��'ׄ ����?��_��(�F?�;��9@Q�|�C/䠒?$�>�<�P[�ڨ����їC��o^�4oY?,�8ѻ7Ku��.��4T���rm��J�4�\�X��CL����|qN�K�v{���пN��h.�疴��LH�U׶in��:��%�m�\[�u�T�Y�^é��9�˽-fs�h�)�n:��={��ͤd��g1׮����s�yeqި#JO��}�y���N�Seβ��{t�[�!!!�5���.���N�t��˒��M'�N��:����uۓ(�қW�T����м��{�Cֹò_���;q^��<R�D���յ�F���jt�x�9��{�s�{h����2�p�R��j�Y���t�i���֟��Ɵ�����R�P��`� ���,�0]$	 >���������}��t�}.��x=ӫ�>��~.c�����<��}������c��]_��>C���O��ߣ���C��\����5� z�D|�P"M����hY<~��x���'���Χ��t�O'�����=�i1�a�iz�����4�-��ϣ�5 ����ǝ?����0���j����k<�/��ϋ��k�CoՇ�����T^����5�$fRR]ː@������+a�V�����.U����z��Iʸ^�اZ��IRm����L(���p�'����n$��+zʾ9U͍��� q���.m����©�E��|�������L$)l"��aN��qjiQ��:;������ε���U�6�q��$�V"�Q��=�c�J�	���3J7]k��B���[���3�CÐ�dtÑ�ÜA��� A<j>��Lc��/���*Ram��J�X�oC�ޢ��`^�'����d"���n�~���"��V�Q7ڀ��n�N3fd6�^k�
�*��^=���L��3co8V���aܩn�fm�ɷ�.8�Rw�eд=�Qg_��h֥��7����zcq��sP���梢��Q9Mu�����b��A�������x#��'��~�������}�0�%:�7���	jEK�[:1�=k:��!̤�8z׿y���&:ˀ�Q�x���9c�`�
(H,��Sy�7<�y��Sk��9r����%��x������yV�}�U��@������N�Ĳ���${b���ΚM�N�ꨓD�Cn3t������rc��|��8٩	���ғz�E���bT��OI�t6w� �x�:��l���̦:�"��i&�6��7=2��^d�B=�����SՊD�e��d�����v6>�j���S�j�5����!��X#	!�W��x�1;�ࡏ& 4ҫ����5�O.�㈰�*��~���}����xRl"l�=��x��B�L�'�ݵ7��J�SD>�aןu`Z{t����5/Lyi�'O;b�9B���z�+^��Hz�w��?�O �\6�ƫ)xWĝ���;
�<l�"�3��T:�R2�y�/Ra����B�t�XS��� ��.�l:��s^9�����)�3}q�>�����[<<��A�(t٥W�0w'KY��V^mwXU1-�Ĵ.�����2��J@󝯜�tK���J�<H�Iv�a����cv:�S�J�g�ܝ:�"�P�آ=��7X��77�K�rt��x���09Y��ZN�K�`�q��
vH�X�wta9�-���@MQ��ρ���8�c��Ƕ)W1�^��Ewֲ�`�|_h;�y�u{T�M<�UL=�;ޣ�yr$�)��i��0Yήڄ�tbV�pt�9x�������rʞ��Z��r%R����M+M^[��e�D$�rt�.�q%�J�l?OM~|�zC�@%���(�B�3�^�������J/���ZȠ����7��s�ф�BI�0�ϧ�C�(�:�g9�֪�C�S$�<<.=�E��r'�B��;����5\	�U�z�E�`h�!��qO���<�S<pE(��p�d4�E#PN�t+��>yu�gG#(��#��GGU��<��₽�%y<$�B�	W����X��\���ny�V3]:��c�@�A�h	:q���Xgk�mESL]�O���9�!a=J�g�<��o��_�0@`u��H`�AAw���1^y>��x^���8đI.�Һ.e?�0�����g[�R�t���g�j�y��n(�'�R��-*�nyJO**�<�g��h���艁�lc�����|����Ӌe�Qs�D���-��7�eM%�����M������ܨ�m�$�s$0��V�d�(cd�wI�i�7��P�x�u�ZF0�
�d�s>/<�ַH71��$�=w��y�˭���Y�m�����hꋟF�Ӥ4�d��$���%�?:o�9M8N%���S����`#�]�6�<h�FS~�Mw;n9,��v�A�[���]X�I�pp�?��W*A������R�A#�A�E�� o��M�v����x����1��nk�m>�>Ǹ�c�\'��w�����w�����I��W�޶����o��|-�ވ16;�ջo��7���U�k��Z��ǫNJ�k.R	J4����7Ͱ��v<Xc��k�����xj����I��Hc�#�+j䗴���կZ���%W���s�_��+��	�%HO0q��<����-��H�b�C\�)G�0�+&��G�YgU���f�j�K4gG�YW\�;V�%V�:��za�Ґ��TF��u��"��k��im�ҷ~�U�3�J2)V�X�4���]�^�3��δ|aL�2#Zh�VYf��%,��k)I�ѭfc��1��Ft��!B������*K+�O�"�M2�� Mc�g�5t�����ҁ�����=����� �FDN��V-�������kI��Ov������=��������_��.�/a��I����[���n���_�o�=O��x^����{�����q6D�E蠢�D	�(�H����
�⮳�կ��ީ��` �Q��E��BoT7~��/����V���� ��K�����)����Ⱥ�?�}�����c>~�]'�ߪ?5E�yƛyG=o��|���b�	�/uH���ٿ���ϧ��}}r��,c��2��1�ȏ{��W����-y��K,aD��,�2�~-r��j�^X��xo�_%������sܿ����s_\�m��7P���D�h=l
�A3��

<g��~/��>���;.�������>޹m�i��Oc��_����q�~O���~�����^Wn7R7q�u��.T���y&;`	UE��Ho�r��}�V�u�!ZY/�$؇�K��?�3D��U�ݽUbf{�]����y0Y��.�o����3W"7�(p;jm��ٝ`�H֑��"���&�C6r���,�@�Y��~@x�\�REB��Ͱ�1�(=������{�/�����s��a�oݯG��=����v?W��ӱ�;��<���{� ۶�h�v �몫w��v�
��?3�D�E��=�=�����_M����d8j���Xm���l�__k'�u��},�]������w���3��~�k�/�e��!0��p1+/y�_c��kUn"����z�_B��}����3$��K�}�B�н��(j�J��Q@�R��B.o�� ��V6AӶ�����ĺZ��|!֐r��}�Y�!.g���>%��i��$z�#-iT!��4
*����kk��B>æ׽�����~g��W��I /����}{?��N��댥{��jL��#]���Ѥ�s���x8 (x���c/�h�#���:�9
���j�R���=꫃y��C�ZZg����AT����6t?e)^%e)�T��m5�u�翗 ~�g���ѯJ�����G�q�A,y�^���|������B��K(��	��� ����sE���)k�fv��)��g!�Ϝ��V�/c�]�T]�٠G�{����:�0J̱��bң��=�2x%�������͠�s�tL�Ճ)B�g>�5�`ԃ�\Y�X��$�ﵞ�1�缡Ř�P�����R��l��ޫa6�w9A�����0�'��oR^*���<Y��3^�f�0��F�x�ut"MB�����^Oh��뽅~-� ��_�5g����p?G�`~���x�?MC�H`��)q�D�{��!Pg�zM��T�C�7B�1*b����mS��$�?xg07��K��:��.7N��I�~��I��m9+	�@ZJ�,Ue�~D� ��	ah�hd���9T�%J�fAI��E�h�Y?AGJ�*�%�A�\��=��UC]?������~��8���q�^�P��4շ�ݚ"()F���_i>	g� ����/�������R�5B5"K9���P���:�C�H̰9#�Z�,,�Ҷ�gE�Wf�*��>��ʂ0��b�x)�Z��⑱�	���2�~�b�q�-�V��2�t�'L ��Y��l�^`��2�/[Yl�hc��M�/�?��W��l��}�!ϑ�����NF���^ʩ�l������Gj����v1��_5��;$H�f��<��(R�F)�e��@��m`�����L��	�%�s��Z=��@�2Jq��}��;����C|�2�K�@4�Az�R���X%a2�X��ԩ�l�;��XÌ#,�f���M����P�3�a�|3�3T��Z��!�Z�}�5�{[�q~ȝ�m�I��(�����_U�*K)P��v��iZ�
̱j74��?0�:;O�(�B�}��c}Ԫޢh�.Nm�F3��"_��<�j�tg=B�8�y�d�F���J�u/O��H�m
�0Ɋ:\���F��?N�8�����|�F�1��b�|��=�N�0��k�!!S�U.�����֊N�h�ˣ�"�[�J��a�҅���q5 _Dh>�Qw��Ү�K���0Q����hsaw�ыZ6{�RЋsQ�^,Bw	L`��b�E�P�^J�$Nv����dGL 01�J�P�RZԘ:����o���͌T��Kss|,Pe�˰���`�QR�-�N~��RiOI�S�*�RB	H�K�(je<[�${"^Su�·�e�(�LL���iE7��ɣ���t�US4�f�h�@��9�2��Q'�Ƞ1$h�Z脇�ș�|�P�.�Ō���y�`sКF3n_�G6�����5 ����Q���~~�Bٰrt�O�<8]7jG=p�X 88�QxǇ��B(��;��V-���0&A���L�[@Q�r���r$"o,�^��$��^zl$�����Ű����V��/Z�fI�j��XZ=��l/B���'���X���8�%�{���̏@�c���-�^2&�]�(Cq�O]-��f'�e`�V�F�m#!�;�:��]�r����.G���s�e�Yɑb��E��Ά�|�-SzU�|��x�9>����	$�@��ok��]KJs��7�*A��d�
�YU�_�0!�$\�L~���g����DD�"[IWF���j�d�����A
'�z�:����W�B�\W�9�!�6q�[ej�A�&��x�]r1��2�3��zg�|e�'3�F���YOfJ�s���(��-9�B�,/��[E(V�gA8���#�]����v�/��(���A�"�p��������i1 ���;w���0���g��)G��`x3�b�.�@lm�|��%�G�O3�i{s5e���T��K�]�ρ��%l��H'���t�hd�g��."ܜ�?���2{X�Og�;���������~��,W}-A M�|N�/�
&��CR�jү��z\�J�#BpB��b�6��b�O��Zΐ6Z)`�$��� �\FR�d ���K.�B��O��s�N���PYg�.�W�B��E�Y(꽰��~��zO	����`u`\YS"64�i͎-cd@R;X�<� ��zV7���m�E'��=�)@^�.�H��'�X4�,YϤ�l5���i~ln��KP\-P'eG��-��k:YUr9�A�	~[�p�3��DДE&����na���"改G�Rْ�^���:�Ut���$�P�m�t���M��1E��E�2A):M��t�#���P��1��n��@�2!H&2�e�>q���`�T��pS3�e��G3o�޺�5�pmIo[���Ǡ�2:�Vst�z9����0~�u3D�o�^��1����R�$����+"Dh5�͂H=���O>� 7�wQ=����֠�Jg���m�%;,f<�h	יQ菭j �AfC1H����.ѿؑg��_
!����' ��=�%�Y:7y��>QT��50�_��x)��|�x]j&R%|I@�whސlY� �>��0��ْN��E(�ЊI�!�e݄̸��[�\f�*.��BN6���
u�zB.xS��@���*M�^y�o]�lէJ	�RE/�����i3���|�!@�"��-�����w��:�EY�$-��i#3j�R��#�I+aF��2|��HH���7=^��*&����r�$�ġ(�!}b���YvKY&,�Ģ"���&����[�r��&�DǦ�a�yM���\^�M "nF���zҲ@,j��=������-x�l\ ��:;��@�b-U�z2��HC$BY�0B�FG���+��ǮO���!QH~.�l�|i3JU �C~)�Q�[If
YF��z�%`h�{�c�8�&"�sP��
"�P *!�ָ�ʥ���������Z#"�k��C��΃I�XPfA%d��"H(��J<D^���=� �#S������/���˜�-_�q�!T(b��p������%��2����\X��7~wN+��L����c��'��D.NDB%Cn���3��}y�O�����f�䤳�q+��Y:�{X��-4<-r���DD�؂B��$\��ܒ��P��؇�w��8��1��,�1^Y��e^�2k P�J�HTD��V��>��hP:�#;���Q|��� hE�g��6�4�DcC�\��P�BG��'���w���=ZY��R'����F8%�-e@?dK�9�_r�ϧ��n���{�%
�U�Yc������T��yQ�i�f@��~���#*��[��4
���hH�>�%��?W�����Q)"8�r���[R� �iG���aTT���W߳��)��UB-�"
�*@_�&R��JB�Z�I^^�Ai�Sx��(\������ȍT���a��TK��ٟ��֋��
�ꃳ�D�(D&���!�aA㰃R��2��X"q�hE�"��O���V ��@��?Àʧ�IB����$�N"e �R�Q�(W<�yB%ٕ���U'���w�/�����$f�2��Jv{��h�'D��W��A(��|���P�T�L"w��ɳ�������wyCy��<Z*Q��\���jl�D�4�{"��q{�8�1d�(�0���Ѳ'M��F��VdDBD�	w{�����6@hH���b�K��g�Ay�fȈ��	���OG�x��K���e7��!0h���.�"Cwְ}b��%r�q�~��?���3����}�:߇�1fE)���Ok]�Z�5$�'`L�� ��Y��@1j��L����.>�O�&O�V���	�-`�x4
� 9�{�j�����M�Dؼ<��uM�еF:�*-6	��Y�96�G������X�W��?b'g�j#���Z2%��h�u�����pg9<���?L�{DB��?6�伞�a*w�9AE7��8}|��?[�-sW���A��=�!L�h��>=�\d^N��=%eD(��0̃��?�Q`
e�%j��IP<�A��6�i7�j�!s�Mt�����=��aQ�W*���U}��jY�.L�,B$��TBL0w�>b��W͚�!D�G/������l�v`��zf&O�É�<;�i�G�w�=���>a(d)Z�&R�MQ��L�4-X�"���'TQ
Ȥ�'�E�q.�{B���ӫA*^I�=S8#Xi:�d�(�#�U@���� �C;<V�R�Wl�����X!��P��~�d�b��\.�TU�A���2yB�R�H\z��|M��ؤ-�\��sCS{t�P�w�ʣ�Ա�t�%e�ъ9J�L�R���UĊM���2`����"I���b�����0y���c!����L��7�ߦ~Sv�O���=���B�!eVA�dR�.m�^����Ş����Q�]b�u�%�: �[��z�I���!T�&U�ʌI�@�_N8����TK*T=�T+-N̆�S@�k���r��U�8�4=%+���EE$�B���+B �V�$�D��'T�ݻbB��S>�g��?�؊���TS%��&�La#*�{�m�!G�EIU�1l&�2���j��Z�d���J�%}��B�˘�TAz�L;���0y'�݆��/$��U�PJ�eĉ梁�Vs�JV��)ZQ
FޝQk
� ���3�¥Q���V[���ְ3�M�GJ�:6�����@��2�ʢ�y^N�K,&,��"���HA����/;�ӳU�[+ʢ#�c��'���B�]�B2(A���N�#!�J46�޻F�eW�<D��W��FC��Sr���Fy��/.l�N&f3ܶD?6Q��Z�ȷ*��qy��T*Y^w���~��=VO|� �P�A�d/�qx���߇	ޏO��.��0��/��~C��Zun��RpY�Br�̉�sm ��B#	�CeBM$�����$�Յt���d��e��3��ʁP!l�V ͫ�"&bQS&��Af `��5��W�^��N���@���p��}���� ǿ�Ƙ�^�;h��X&��`" �Z���KKYD���w\�{���e{��_�ױt���ޙ3&ȱ�Z;n�-H��54u�_���
�>�\�}C�jD�'И)�D�|��0D�dl�z0F3h�&9��zg�o�Ӿh{�$vV�)Hj���{MC
�UY<VJQA9Z�LP��c����ǟc��WǢ�d&�t������,R�dr�)�L��]6@�=�G��Esv�?}�8�{V�$��U.7�$��L6��~�,F�'��bu�����P���j0��vD��C_k�"�r�����X�	(�k 
������C0��?y�oB��U��4�U���]L�]�U^�|H�E��>z?'�	)����7��Ĵ���� 6xg�h����Ut���&�C�1a��H�\R�6z"�E�$�=2�1@������'�Aʳ�%�\B����h�$�Ѳ�&D�ԡ2�Bՙ#��s�M�Jd����}D_��u^����e���#J��9hٴ�*��ӨU��U��������L'A",���̮����Bt�5�T��f���?		S�B��:zYC<��+W��*q���]�|�����+4���<:Β�Yt�׍)Y�,���6�Ed��#�oAÇ8�Q��D�_N�R[U�J�;
�T�J�������R�I1����i^΍�+T��v�)��f5!�=&���~Eг햽�����W#Q��H��(d\�|�M��Aa���p�^�Y��"��ա���ZR1���2�62/�r�$��]_�{�S�i�A1coY	%�2�'��Na��KX���$��mB�1�D��wR�L�TRxhE���r�i�	������=g��(�ZH�.h�;gP���1��= b:�,����߇����{��W�8��"8����4�Je�r�����a�g��� ��3ʚ�
&Sd�V�!�+;	�թ�XJ/�ؾ�㘊ho��p
 ����K��O�;Jzj0׊F�����_���|����[�ʐ�2�j&���<řP�d�G(e�"��"֢�~���^A|I�<�9�y�֨�)�Ң���6 D��(���Y�P~�Q�Q?�4��x����M�8]�h(��<�Ȳʔsql����QeTT�*�iN�������-G��	�U���s��gY�� ���[�2�2�}�C+��Mp�%·S���M)AYDQ��-mV�����e�Q��5�_4[��
�xAJ��̅�0rE�Vr_�����L�fK�`)�F	��d�GfV`�d�޺��e��DάJ@A��V�/}N�x�,����d	�r| �k,�����+���F(a�F'{�ZtSf"!ḣ�^Mx1����,3�.���/dX�C��l:�(��
0� �7G���+������]��0�Z��>���ϭ�*��(��M`�m��^o�E���Q��f8h�Tj�E����yT>%`U�
]#�uȵBƊ�\%�a������V��J|���@��%��
UR.��?�n��FYlT�q��2���)��n�'�l��Ꚏ�V ��J(�5���[��3EZ"�e����+�wɵ�v%�I�A����FE�}�K�_�;���b�>�}f�(�d�*ơ�j���C�4'(�	JX6��G����Z�ޢ��R�A,�����N��%ڨ	>��/Q�����:�%]c^/���H�������Dl؜�R6G��AJ���}c<�A涰(�'����DI!BMJ-��.Hv��D⠛�6I^/�U0g	,��`K<$�/�b��tV��fa �FfbE�aJ�o_\�	O;6�tY2C �B_z�_�x�9X}3ֈ펀Aڔ�2*������o�<
��N�tv�D�I�e��BV�V�i��)�oq|�&RN�A�@�F곭M#5{I��-V��:.)lgvj��])�e\�!%�9]qY��A�\b���X��$�;3�H�v%���wQ?�V�y���G��.�g��/;��g��yG7���{�:��Q�J0�C��eKi\b�3�Z�[�(�ai&-Qf����X��'�d�J�������m��2���K���!�#L�di�������s �����+�=�;bh�y}�m*�D"QҋA��&��1{܋Y,Rf�����C�=��Q��]�h*\�P���V;�[��R`�Z=AET�ڢM����)cj)�	�(A.>�6�mƗ�"�i�_�DEj�+o��@�"hՁRc�I�qm���l-��{��*b��K�ZPJ�fj���Q3�@��e���P�ikK͡�1=�H��V}�8�~���ܥcEz�X�E�
�7�e����"Y-C9����ym��0�r�okS'e&�B���ל����N�4�Z��(m��%���F���oK�2�����(e�U%���$�4�i�_�Dy��2���_!H��6.R��͎��혽��)�.�.#r��l�!Y���W:���*�(pg�|Zc2/�$��bjh�6J�C�D�H��-SMk��ԍ��B�F�EvS�F�v���b�g�I��\���4(A\�lF27�Pb8���}�~�^.��D����!9��G�`R��nD"5�,��Y^3:햰U���D�DҢ��2���R�,X�f�b����6-�;�NO��X�����h�xY��ཫT��tY�f�`�5E,'�V5��D՟��Yg�GL���R8H@b�m�r2����X�Q%)~��3�������K��?�1Ӯ�D��y�Ct@��%�,��6K�˩���4��F��%c~r�R��#"�$P�^�1f0��p�y�"mc�0\
*�ɖ���	DH	
��J�zT�;��v��a��v ���R�Rh��Q�c�LI�,	�*��W�s�x��mI	����
����J��䛌�
�FL\�I.�'f�����W!]"�(�b�/����/���ݤ�
� ���$�u�.�n(����(E�3x}$�hg��,A�D�Z&R�5L�V¤��:�A0{��j��Y?_z��5wm4�t�@��U�B�A���?o��k��<>#�� ��"�1r�J��_z��æ�`��B�$(�1iT��Ƹ�h� ]��o��Z�?d@l
!q�E6~	�Ң`�K��rR�Z�{
v}-F��b��["���iZ5A(�aԉ�,��o"�:U��u�^n��
�)�9��iV|�]I*�^�IR�.'�2�?]F	�L�&٠d�=����I�@�R�`PɑF^�Ҍ�-v�)k����:4�F��&�	M�N�<�Ŗ���UB
�� E��u�n9��� (K:Ņ��3B�Ie~Qu���ψ+Q5N(�1��\־��I6C[%Y?Qm�e+V��]��7(..T�K��R;�Nn����wF�-Z��tD0+n��A{�^AK�8ƙPC=��DT�.#Mc0dH�JN���˯l,&2T.R��j�Jܮy>x�\R�s:!���q��`J�.����C!��Ԝr���Q�"@���M+T�hĸ�U\��쫼��}ЊV�
	����/�!����1U���IJCk�
$D�A�Zh�XB=��!R]bD�$]0&���Y�bTz��.*
�1�4���|��IǻQQ���2�@��F���T%���jj�1pp�K#�֛�2��U��j���ީ$���u=9sF7.bf�=�zxݲ$���]��;;
��b����(&D� g�	E��9�b�	�OF�%Ă�v��]2�~��kЀĂꪲ�A��m��L �)5�}{�2�ȍ���|$ >_4�29u�	�KaZZp��aU��'m�(�u qD��\(�[o�j\I0!
��ؘ��:�K�	H�nC*@�_����##��~���a�0I?{�FQd�L#"��C���#���Y��h��8��k�H2������F��"q�TU5�&H��b(^�!X,�_�Bã8��,&ԓ
J �H�v��Ŝ�t��y�&>?9r��+���Q��),���M�K�)q�-��@|W�]����F�怆�O\zR�,@�@� �0Jg��n��Ɓ��3� �pQpUR�f��{!�f�V`�W��#-��ƠP�������Q4��!o<�3aEtT4�5�N�Ir�@h"X�����=����Vј!;�A?�_�a	ù,"A(��ǆW�Y_1�������7��p���������xԦ��4i.3���I%@�QȄ*�0�X@ᒴ��ֿ��ղ���D�F#��ő~�9�:�y_#����q�T �h4>=#P���XIgO��ė�q��ŬI~����%�| w;�h���M%=P����@Ֆ�w
�?�L���X�G��N$���D'&LPY�_$G�*�D��[жS��
�!PA$Q�?	?ԆR����]��lt��o�|ן���`��7>�1|>�O'0۔�S���,�E%��d�ބ��I�
q��E{D�����H��`2��x����{�@w�#�`m��v~��!M�FZ ��Lː�M|}��X��:(3�(��c�O�i�rBP��iגЉ!�p�+�h�W1�`�1V����E��]����Լ�ȅM�G�GG$�s�*�.Q�bL�,"�_~� ��g�O�&ww���jG�ȏfB�̅�ܭ���:Qg$DD13��D1I&�Ļ
������y����TNT.n#����~�l���~���՗q���B	����R��
�{�.���L�5�G�|�|7���4}���˄�*]R��B�o�ŠF'%{��?Q�J�9����5D5�hD��ց��$x�Ye#��, B�U�j���0����3�W�+�>����x�����������h?�dp���a�P���<�	��|��E�ҷp�-X=���@���c��z��By:���ε�h���F
Q�R���L
������~SWOҝ2z�Z�����b�
��Қ�f	0�k�>�	~���z3���4}���1��	"��Q�
�����A�*�ҝ�"���376�D��T�+�X^����*J��}`�V��B&+�~�s��6��)� ȅe��m�ʨ��
�<�??�s}��k�d�(6G��N'w�#ܵ���vD0Df�z��<|S���1?o/c"X�D���@��Ţ`�'��O6N���7D�
��\ty�&��04��;Z��X"��$DML�.yD��]~����g�=�8�G�����:���N���0��I6F�+��x�M0����4~q~��zR�J��Γr�%R�w�3t��B̚A.y�*�q����D�|CC0��}a�VҲ+;]�^E�g���T�oJʡ��+׾���T�fiv�����+�H�5D���P��Z�J��ٛ�*fX�0eD����h�����=)	�܂�L��_(Y��^ �3R��(��Z�������QP�aR��&��_4gބD�FQ=T���՞>`�����P�}��&wvC#�O�y�����sM��
�=��Q󔔹�B�@E�f
 �%�[����##<�+X �C�1DD0j�sj�+��^�S/�O�����͈>\��7���#52���<�9"��G��4{����2�5�Z ����.j¸&W���A�Q���)�	Dz�(�م�]��]VL^����l�+��{ڮ�`�,Te:2;�؄��L(rg���X�+}P&b-�uAz�=��(7���n,��1Q-�M�YX�JetѫsS���m�����6��{�zRQC�2���~mP�-���LǎD��~��3��CN�I����*�8�����A���Ｘ{��D�diw�J�����/�0�Ӿ��~=�֭>tc��!��m ��>A�ȏ$a����K�_��FY�C\Ϡ�X�}D�~ѯ?��? �1��5�2DM�z���O��w�ɝց�b��V��

�x���*�.(������4|K|~jL�a��A��V�LIC�dD����sxLAig�38�SG�]C�+�$�� 5OޏiQ���/��^�S�%{��~,_���||��~��@�-l��~C��8g7�Xf=F-�5�qu��I�~hh}�}���/���c�a��?�w�#A0="�p(2��H4Qd�E��=̪C���1Z��R��7����)�c�d}w�z�}�Ή^��LBp�K�f6������?AK��24dYM� DՒoW�1�?ccF���vc�7�.�c�_�g�P6"���l�N0D%N��K7��V�dB`�����bǿh��@��J3)+Ar�󟟶������>þ��v{1�B�l��|a*尶O�~�S�^
�U��RL�����(���|���
��UZw��2��=$Lq���U�T_��Jb[Bb)��#6�]Y`�¾�#�%je�ж�|-��kDt2_����Ǉ��ۙ޲��ι���d�f&+!$gУ-e`��&�K �EB:q�6��i�AK���.o��M�9n�Lڂ�4"T`U�T-�gjZ�X�\F��ݐ�R�V�e��X�au#�_x\�L�9ʓ���j�%��y����p��	���)j�3{����	L���Cb���!����g8{9�s���g�$$�V�m].@T$���hr���0J���  �P��F�T@H�D"�"֖�J՚��Z�����C#!! d`�"��̪(1v����
(<��˄�DD��ѭ�"�����e��D�E\M�E�#�����?�����_��_e�_�_�����~��r��P�
���O����$:^��o������{H_g��g�����T�ɐ�ȼ�����,i�K���ۯ���Q#��r�a|�!'����GueD�'�{|�t�6�Q?��wf%�P��7�z��.l�{Xݯ�_���(�.�!���)$<��f�,J�	�0�R��\�����o�5���K���8�Q�ū����[z�7=������M0U��B*EB(@��I�	dT�K(��۝�)�O�@_����5j5uko&��dU
�b�u}�z����Pj�H��B �W�=�G������dG-"�N��B,AA�=㉽DƸ �V�:F�.��9�N�VA/AH�LҎ[��۷�k�������,W5J�0�H��Я���7�|�����}w�/����O������?��US�\6~����=~���|��W�����q_����t�d?�?ܠ����ϻ0?�!���g�����Hj?�=��cW��u(�Ł��?��_�������&�f����Fѯ��oru�6ʓ���b$ ,�@	��	�=�]RDK� ��߸}����j� �D���fֵ�*\�g9�([�S����z�o}V 9� @����׫=��������������>��g{~���}6L�/�迤7��G�����������>(�������.���vs�S�H������m}����?�|����b��h+����� �G*r�U�'1�3i����h���v�zV�W�����?ޗ�2C{���*�� n�#�f8�[i����$�C��9���U�N����}[V�����N�6c��R��[xO<��p��yֳ�Eh�Òbr8i +�u#�I� & �  '�8�Q���~�g��C��	�|bY��}��i;�%�>������_˺p�m�������qw~�E�~��,o�+���RQ4����*�ӿ}p�JVQ9�aT�D��)����oM%�W?~����TAH|�-���v��#�����y�>��:�D�ʿ��:��"�̀����۝��VO���1}�I�����6��0�6� <oမ�6%$y�����hU��%�q�\@2O�G�"JYꉆ�5�.�FщD&I���wZt�iE+e���ěrQ�����.�L����%-�@�/˘>x#ԇ���B m��︯��sV�����n�4�
#��@0
EX	Q�0{0!�/o,C~��m�M4Po$v��
�x�0�~�9��h�����;P��p8_?��������6T ȡ��YROVW�H�[��C��?��v_�����cj(�����H�|��̓��"\�3�.���oO_�~e�����[���o��*1 �
e�G������J|� =^���;m��ݜ��oǪ)�fx��K����S��7��A�˃{!�N�>���t���ߧ�lׂ �XD8iO�J85O��<�u)p�!��W��W�������Y���}7?o��s>'��#�9k�'�h_�熯	�t:��Y�g!��rF��r=V4�O�og�2�=��z>�y���h��K�]��:�d@>Z��G���'�9?��ߒ�����%����(�"O]�?������.=9D^��<��ox�����l��7�4��x=�}ƨ	�'�x��������>wJ���]:���W��8*�FbP��|�x��o�?��vA�{�����������(�����}�L��!������5����{m��Eh��j5�X#ih-����Ŋ����bM�X�lF��E�!1��Qlh�Tl�ّ��&a�Ƥ�*1��5��F��h�1lDRlRcm��j5&�_�����{��_�Rڧ��Pzj�<U��;��N�w:�3v�(НK�?��N�[|����"C+qcϹT�q��ө����I��dlHOl�EDr曠��S�CH�o�Z�.jC5�",X�0V�5KW9\�]��wv�\����Ƌ$�IT)�L�֐�w]rݻ��q�v�\��P��N�k���g]u�m����Z���(�b���-�F6F-��Q���Ab(d� ��4VH4a*ekk���w~��^W;�W*�?�?�)�88i*̦U+
2Q$�Z@�%dgNe뼼t�ܺt�M�],r둅!�j�5�� ��@ �B�j�'��E����������D[�o���������"�!�dݭڤ��K��8 �wwM��m�S!	���BS*�[�km����a�$в�V�Mem��bQ����T�)��*��E@D#�%8P=���ږ�V�Z��|���7~9�|��2�B��Bh����.��^9��^-�
�@W12�a��2�ac�I"�\��떫֦�{v�u�I Jݻ]ݗuC�]!@!���H�bH�\qq�G]�4RdJ,D��2�mkj۩L�%)�6�mz����u�g4�]κ;�1$�:��E�����-��n�b�.
.�dQ"2%θ�bs�M�ut�:�ڶ�okמ��k�ru.I�s�r]��9W9��s�W.��Z�u�p���(;��'s�ɸ�rJ�ws��u�9�3d�щ�i��X�:u�q΋�P�����Ub �0`��Θ�w�9s��g]r.���;�w��D��� �
t�JT�7�V�7��P���B�G��O����lT��Y
�-�0���%��A����і�	1�*.+ ���+)a�!X�Q�2�[�����[mL�B�X�BV;+�nIc7]6.+# U�Q�m�U��[X@$\(���!K)wn���X�D�*�-hd0��H��D*��ڤ
ī�A�����Y.B��$Q�d&��mr֍�$�L�Ӝ �"�"��׊��q�&,iMk�k�>�eZ����im�`�%H_��J3����m�H �SADT!��L*�s��1v\e�L����K�(�x#z���p�I-.�ThG.���ӷ��w˙D�EF�IRUm�l>L���o�f���/����|%�%��n��et޻�Ǯk�'Jo;��՟������D��>��'����1��Nd��SH�Ȭ�H�y�z\���-�ny�PD%[-lf��P�I7!L<�Q8�L�H�������,�v�͖rJ��\���c,2��v���׋	:I�B\��ȳ�����'nR.�l�Fqr`���0�Y��ŝ��w��٧�����-�e��R�lUa=����Ge Tj\2L��m�2'T �ʘ�%$�DKF��%УIi2E1���&<����vn��V���+���YFT��D��LeV;yWh��FL�s1Qyat��2\�3&�\dd̬�M�/31�2Ԧ\LF7�kⶋ֔��_�p��ZɛH��\T��t�$ƘLy*�+6���C%T*!QI$��Y�ʂ��/� ��!yg�3���U�!	#�,���!��i ��-0<����v��^*��E�ͼ*�v\sn�l�{h�K�R��"�*%�ǆfJ/%�*!�L�Z��&(Y�#PnS*9P_E��%��V��b����: Q.���c���`˅Ʉ2^�͐��Jh!
���l�9�RѸ�,�Ht7t�]9�A�������2�.te�:0� d��:(b�q�gc�B���Lp$�S�{vdL͓g͛2x���W�>��Λ=��@��\����>�6B�������;=�>>�5�&��x	O���R?9�Mٓ��8�:��Jn�>��'�I��|33��P�lB�X˖L��/��_2`�0�v̸d�I%�g�pnV�$�9�3s!���mٛ&�r�1�<c����)v0�c�gG3�6o�=��gO�[��RIf��`�q���,Ӊ&�de��g�,��:}�s�Nm���p�y�ˌ0�HϮ�n��0��繙W��$��f}�n�q� d�vZ`;8� ��`�L2���B��P��2�dV�5&9
�*!u��ff@� +Wa ��	@8EQ�W	�:��̅����x�٥"}�>�S	b�,�EM$};��N���Z�RJ�T�%���V0H��ia�[�IhF.�V�QR�n[nKS#�1�6%��~�O2I�C����p ��{@�-B7e��Kayp[[6 a�c��C'Xx��_���>���r9������H��:0�,����cL�屗œ��@��[ay2(�.HP��Z*�`��Ȁ�f^{��f��H�ڶ��}�n�ۂj�f�jR`A�/^AM�vZnӕ@$ @T1U Pp$V��|ɳX�� ��n�
R��Tm^׶P���A�]8�]��s����[�Nw8����߽�m�{���ѱl[�\�ڍ�+��r������������}������� ]k���o�xL�4,�#m꼿����m�Y��ĩ1���
"�~_����7�]�׳E{*U�����j6(�F嫘��-�\شcZ�ă !��� �bu-+i��e�el�nm�����n�_�~c��j�����$�H�	(ɸ*+r��oP΀2[��n[X���nj4V-�
�� 
��@f4�@���I��C<KI�|x��x����������e�`�A�1fJ�22��F�4A�M$	1�sBw\�Pf!�׿Lh{`,�T�0�-�oK�:N��8x H�"1�W�b��/�)���OӭR�6�P��A���e�����۹\KH	��͠����Y7��HM���� �S�����������	�����O��DT3�sݞ/��D���\�dZфYH{�v|7��Lx�������r���J?����O�`�mg��8F�?�0������<�2*�"�*���f��'�N�$HP�<�	��٠b[�o������1���t�[��sq5t�l�K�H�߆��C]�9�^~�!*\� ��r��_{�
���w���/CL����Hî�e$�� ,hJx�����3eG:�?j-u��X]���91@� dU��|}b�=
>�����+�a� ��3��C!���1/!��@�!��������Q�̖��f�̒���Al����Kxv/�d|d���E@�tB1	�����C��, :_q��)!'`���Q�h��maK$?�F�nSe"SQ�y^�b�1r�$"�U|/en%�5gʗ�ܦ��0�'���Ͼ� I>	�� NX��퟉�	�S�6�Z^��<��H�a�+�EɎ�q��(�Gg��|>S���+Θ�ޡNS�ZR�O �C:d����N� 
��d	ܡ��= ��x�g�4����ԡ�/��璖K��y{y�&z��/w�'�� x��	�`VED$dP$'�ZyxqTt�Y�����{N#�hz���q����T_��o�}��O�a�Qn��3�LK��]?��������������?�m�߿�����O���_K�����ɠd�/���|}=?I+�~\[�_U��ߴ/���?���{�*^����߸:}�8~�����G�W�����k�w/���|6����2z��;~�����\>_�������O���?����_��^��_�oGS�=mK�?��ó��[�S�H_����Rt��We��)���)�� VP*;���/���������0���hiO��t���z|���y9�����=o��8Mg��5K���j����r��7'J�W>_�~	��E�K5����{/C�j�0����W�i�h�)�5�*��ɸ¿�=�ă7���|�?"$=����U4���<�l���L?�޵��%�!�I���oO ���b\�Ϥ���c��d���Ғ�Z_��Yq]��B�ݡߟ.=�	g�G�'��Ӳ�ƌ^~��rT%6���(���������ê�(��n\��T��/�S��$ԓ'��9��d~愎�))�Ř/�y�d�$h�ns��꾈xA���������z�N%>��9d5��{�vs��-u��/�x�|L��J�7���W����?H���i���i��}f�~���>��v��]�_�Ƕ�o��A5�vɼ��m"���*��&�E�)0?�N�,A��R ����_�` �t�$�y�Nb��	��; �p:�����x���W���n��q^�/z��'�ƠXC�:Y�z��,�W���7 h�y�y��������RDFD@���D�
� (���vΕU[����=)@�_ck�w�� �bhD)���x��QS�=\��r[�ԙmλ�Z���=���޿(lq2Q�é7A(��҉" �|}�l�!@�U!�i=��P��p�QK�������=G����h�<�)*�~nϏ���q�j�Q� ?U���&Ъ�5_��]��t۾]�4i�$�'�L�Uj� w=��q! BEB@dDN����
�J�P��^�l��ENW�������2FDx��p0�.��ͯ�և��;��m�W���nn���������|���'}�sg��a�/���vM\�x��/�37�i ��w�*�74�ƥ�]�Ӈ#����};�y�x?o����Y�Ǐ7����ܩ���+{��>��ߌ�s�vL��hj����-r��������g�_�����~�����o��g���W�^���~�W���W�\��<u7�}�+�\G�
��U�}�ߪg����K�~��*,���AD��G�}��� ml`�� 3�_����!P�1���������m����8���p�0�5��/'D�2��̀�7�[�G�3�4��25�cJ�/�=Rg�9��. t����DEY��f�Ӳl��Z-�a�ݴ�{HsUʲUPTd
Oe]����7�,��`�RD�G�#9X!���E���E�C��j�l��d!$l�{�q���_��V�Kܲ25�������VQ1XS[W+kcj�Ko����|�$F1����e��uE��h=�r4?\;j9�5���W�%ηT@҉����c޺�v�o�PtJ��*�]���Q�*�j)-��"�`�L$@�"�S�X�$U�=����ð+�d ��`���"#B)&i)(�☪a���aFB�5�R$*�Hڪ1%�E�
��lW!���$�	�'v}@ƭ��[V���Q���"M{hZ�j�o2�]tP��0�A)�ԝKe����m�E_�����F�x�Z f A=rADq L@�D�8�ƀ��(3��"F�$�4b$�BL�,����[�T�B"D@" �A�p1"܈bB(0
�g ��tzL��e��}Z�Z�	��u�����ީ9o�2�v�=�)�������=�ޞ%��F0	�J��P���@�D\�Ā������E�R1UV�07�Qnq� :p�c����fM��9s�VںUV_iuo�����W������I�H�-X2[)lJ��b}��eĨHBBM��V�⯛��dHͣP/��B��} (���5ț8�=����/W&@vq���k`
%'&���n^�8�����4P��=��M�B�3����\�Eƚ	�@)6#!7���4dFBBA�$�E�IZ�����oo�*���"u�\e(�: �!�봂�\���ȫ����1�&����LRd�9�L�$��"d��e��ۥ��d$�)$�I�"���F�f��hT. |z��8�(�)���.��qn>� d�n������	P�&��t}Qӱ�x�%4��)�Gj\�DQ/%r
��"*��X��K	�ɚ��%�U�j�K���;�
ԒGU1P�U@ؔ4�AVEO�`����HA��҈�@o��7��)��a��@{tW0PTB@D&����7SM�Wa�p�-b�ʾ�Ǌ�(׍��-ߊ�����B�E�sv����
�
�"
��D�D�ȃ@\o�p
��Q T4bn��"�=6vu8�2�c��ȍ�$b"����p����D�A���o�9`Y]�4i��a�PI4Wը��ZT�$L�d�hQ�s��4�5C:2�,E  ��ȃ�	� �l�&�f g��8���@L�fr�k������mʹs�75t�k�����;߄�T��ZHKRS7� j�2��M��I���AM�h�����|�@��uٹ�ﭯ�������3�P9H�m��m`A��Ԉ|��&xf|܃����Y �B$!H�2�gQ@ H�'	�zLI�熺�B����UIDY-E,��-aD�dm�X����$��I�)�vm��G-;�9�4�R%tѥ�4��X9��\�.0��)��wvI\���.e�F���W.�)Xر&�b�-�5�Ӯ�G];w7c�"�I0���H��&CB�o�U�)����4�E��$sw�|���C�82�C@��R
�b �B�R ADs��2RA�F�7��I%��U2�P�K�Fp�� �K�WR �i�
nh������0w@5+��1|x`/MJ��p/�@Խ�1�(cA��2+�[�T*�.a��&�"�.~���7���_+���w��_����u�}L5}��ݣ̭�ů��0d?o�����������'~%��쵷�8ߜ�I~̬���ب�_�FPF!���0L��x`� �Kև����x�{&'�f&IT����T]�I
�Ԫ�@O�I��I�	ə��,�Np�|�W���3a��d�y������g�o �ԣy�>���K?�@H�YԸ$�J�27���XCF����C��١1C�[HQDW����1YU��%8-?�4�Փ��E�)�U���^���+��"�cF����5��ζ�ӻ	]GPWT��}�S:Yz��W5�S�9r[��,�t(D���d����Bz�0�⩩$#TTd$��IP��~���O�x <���4��ܲl��v}-�������L�OO���ϥ�rJ������?W�b�;������=�	��6`���>̰*�$K���)>���h��U��R�o��R�hZy�A � �$#(Ȧ�%	��In��lpn;(������g	z�"��
��K�|o��mg�ڭ�o�U����U��ߊحX�鄱/���]|���U�`���{w=^�<߈��<����*
~���,���I���S�M���_�����Q��^��0��~C���Ǯ�՛�H�T$D��1���xWq܁,��Uݲ����#����sP�@�b��7�f��OeD��B�hs��`���b������˿���n��Ӽ�}f?k��̼��~w���{L�쾂���ߴ��F�%��-��8�V���O��;���������djJ�Pr�,���Q��,R��?�p��T��� �r���U�^Q�� �x8��<��j�:=	�7Ј�`Y�D�_��;c�Ip�h?��_��������G쾯����/���]�ÄP_p��}1������g���>���~�t�������	���P�
E�>�a���G���5�>@���|E1)4�#��)̑��I�Q�I0Z��HCz�i؆0�)��l���cz|�������j�pc"���5���~�ځN���^�	q8*�¯�!������A��gi1]&O0�r�����&���/-�,���M��~t�c�!��P��\�_���8�)���Э�?w�lt|?����Q�s�N�"oI瘷�pW��E>G/�Df��9$��$�h�}��=�Il�X$dI VB���/��=��?ã�/�������i��u&�4�@`��n_.\�)a��(�:��$$.SR�Ѽ��6V)x�0�U�bUABC�)�Er�� �`��"���{H,�H�.K	���0���(bP��ׅ��   iL�L�G���IB�P�M�@�і��EE�G��P�K �@,ѦEO���g"<�
�"�f'�J5(: � �``���
�b�������1e�H
��0� v�%�W������}K?:�Z�������r�6�p) �A@�z��ѭ��Ճ��m�$�H�	 	�T�AUK��.+s��f$����0܃�K������f��rv�˱x���~����>�oc�@2~w����0���#���ʲ@>�/��P�p��Sۥ�������3k����tp�r~YQ�Y�,���k$���1�+᜺���b�9�U���]"T�������#�%�6!���G'
�=Cy,{��B,##d�����x1]|������?/� �(�����������}��o_�/�Ȥh��ē����G�_��!�;�Ur������އ<�(��DP�,Q 
%���� �
d������'�O�B���=���ȁ��G��X�
-X��,���*b�i1gj��?��p���T��k&;Np	ǂ�d04Q��`��H��R @Q`qR)�uJ��\
� �â �5�Aӏ�?^���5	�@<&Y�A��W]�xx��*V��e���n"�B��b�z�M	�7b��%J�@԰C�%�d��cF�� �L�tCmK�+ �96� �5��P~>���. 珤<iu�@P�@��f��*�,Dli�K�ݎ;R=�.H�?(�'�8i �j|�D"��fV�q+ze ��=���F盛UdQPs�(]��`���y?������"}����?�`	� 1���\��O!x:�چ�	��U�v�jA]�28	���(��#d�m�%���ʺ$D�ֶ�h	G�C��w�xț���+��{���A_�m�e� ��]!����@$;�1�����Ͷ��:�G�(őT���l��çq�";^�.%8���������v_��}��<;��"�2
缑��|~����>��)�{u9r~y�'�}9�)��9r��>Y���yY�����<o�8��ՇrHHLYlc���\�G'���O+��v��[z�L!}���)S)Pr�(ȈB �=��'���/�K�d{c�|3�詰���~�w��䷯9㥹�G��W-���i��~^�3��d��K�ͻ��5�;��q�p�~c@�LAư��������v���Y$�F�z���_��f��'f8��.�'��
�:3e���x.�D���ݶ�k�$$�͓Y��1��!��~�a\�*2  Ct�>iƝO]��Oq`�q�,�R'f��1pw� �1�x���d�o B�x@�f���zث�*� 2
#�|���$��'��S���$���瑭o�~�a䣐G���ђ���_������>��<�:�x;O0��y��WddU@Bn�\��}������2}���~m�TjI�i		�O���r����p��M�����������ZO�l?��ې�]�(���� � ��=ą��d���<�� OѬK�ك�n$��p6��d>?\Hq���~p�{��d�����-?c�xBHX8�.J� `�@�V\
z�<_���c�>��� ��s��= {�7��<�E?��<���X��@�k������1�$jURf�(9 �����[�І�v�^	����=@����%�#�ʟ�����Є���|���$"Ke��>Y�nPq@RAAd@	�y�FBA��}N�PU~'p��ɑq e�o ~���m�����b���$��~��C�`)���e??�=}W�$`�Ȩ���M�w��n��=�1!,w^(V��>�,�����$E�t����H�r�dDFAY�:k}��ZT/bq��	5���Y*~��tq����r�����=8�;�2���쀦�@�����"H*> Ｈv�Ph�ޒb��?�h�#�H���q/�bp��#t# A� d�;����[���GM��ۼ
��e=O���;��T���C��szHA�GŁ���;�Q��0����4�/p��~�/Y��.��y}����w</��?����G��_GE�u�7��_��	�p<���7oM�����g�{'7��9c���^�?C�{�G��g��=��}��w���{����7���NW���h*�^��y��������Ϙ���-�D5��֯�ݴW�m�����(��0���"`?thn#9ea�$���G�[�(� �Noh[)r}����I��a���ğ�j=
��c�{`,�c$zP�InFl��P��R�c��ȋ�'>}c����k��{��}1�y?��lb�
 �O���#$�,!����Rcd�Mn�d"��T�����IK��/���P�w-�a��#���\/`E�|
� �,@.��(��͛��!a�������or�i����Pz�H�����P@~���`�@��c��1 ���_a�?�����o_�;'��?�������~��ۿU����H�*?��e���9\��	�����'�)C�"3�,���Z)�|�#�/�e�YAT�m?��XG?��
={��-*R̄���v^^@����:x]�J��C�{��W����{�R���Ed@�#��ߘ����=�퐖1 �=s�,y���px�N$:�yڶ|�(4�T���"������ ��$�8�'*0o"��珤��^D�������t�	���l�|
D�?����
k�'�ڿ}����-�ߊ�����^R�2c�}�?Wzh8
t���.f���!7��[fP}y9�4�c�;]6/k-_ y�����G�N�)���m�2HxT��"f�B��q��Q�>�K�C��48A���
D�^�o��C���5��/uԾ�,9��zӇ.:�bE�Y�8��z��/�k~9.N��� *aC�<�õ�Ѱ�; Q�x���IL��uLƞ��������O�@��Hz�A`>�T'���n�a����&!G݅'U�}�[r뗲�Ɖ��|q��B�H��S�iwC�-"\�`���T��	 G����	z���E3��M̂k���B�
 z]��$%ǎ�e	�� ��#��'�<�&$`E�0�� ��"�EU0���c�5�p�0~�GvO�4v�LX�.����b�^@pM�TJH �]���c�I#9g"�=TJ"��0� � `�*�H�b��$@��<�s>�/�_��o�R����
F*2m���K��ٸYq����L�0�������w}����e��*c����LЄy�'2�@DE��)�`��6�ꖿ>�Vɪ+�iAI "@"�H�����.���;p��Y�5 ΂� �,�0�� ���`���rP˗�����J�*J�U~�~�E��q��U���赫ݧ����T߾�G�ںnӠ ����]�bZ�//��\1jKP$��D���ӥ�t�uUA'G�m�xA�n�Ɣ���V~��������?c��FW�7��Ƀ�x?��0���$�'� �
J����mǹ~R*��pYU7��[O��%b�m�`c��4i��Þ"�**Σa�#���=�q����I�9��uo�{�������rpk�,ɨ�A\��{,�G�E�<AJ��������P�U˗����\W����&B�yD���;S_``�ɓ%d������z��6Nf
@��K-f�kJ�Tե���E�D�H)#b�88����<�
��cA�����Z���9�����#�0��"��2�� ��0��*��La.['�*���VoX,eIF$SCo��_����Kb0�+e3"��d���2��F�?+�*���'�8�Z+�/��4�`Hb����X�!���TY�&�4��o��-�3��s�O���h��k���hB�C	4��������Q.��٫�2Q(#�^V��%�� �" G��I�7&w���hg�FrO�����_��)� �|f���7L4!������f�dc{i'�iw�5~��t���<m^v��q�K)��)a�9\����1�J���6ь3�W[R��u}��k��T�9�Hk7�.I�x���Vօ-"������T85�Z�N���5T��9f�KH�B���p�2�r���B���{���կ0�iѲH���j�6&{-v�e)�o[�1���1�6�(f��a��L���*����]%��X@�f�Z��ͬY�;�g{���&��s�U!!&�����?� ��NY?��i���;U���4�K2�4���K<�[���ߝwF��e�O[pڭ!xi�BO�:��Lr_��2�|5�c�Q�i<^���W�/^Z��oC�ិ�|��6�o��L��8zόWhR# �[��<�L�t��ߞb���,��v�W46�C��u��{æ�k����$u��~g���F��+g�u�C#&iDHg<n���'ia��;�9���$�����u�~qy�o	;?���qڹҔ�P��a��F{����
�
��
m��Z�Ϧp\���r��[?;�B�Y�+��we����}p�k��e�e���6��L���2*�@�UPAA��EP$PRAPEU"�*���i���b�i���c��M���G]����hnt��\�۶5h�~�m��k�ݻT���4���ᴕ��^Gd8�.����ۗ������w��+)�e>g�����.����>3���	m�z�T��}�.b���5N���D=w{�P���q~4�)sڝ2�!m�Y�Κ�;�4;�G�ڭ�=r|:v�A�`��M��]��Y��׮�snz��.c�ӱ�IZ��Ꙟ������9���b|%�	��nئH����g�]���1&�z�^��iu�G������w����7��:ϊ�{ˮ,��	�}����.e��p�f�7\�e[S��;k4��3�X,uh��{�ߑ|��]_�Jq�YL&8��zQ���f�3��jr�Ǧ�d�K���~�Y��GVE�0��Q��_��b�,8�� D1�6�FB��Hd��D�h�3�
��)*�V"R� A+eZ[KT����6�m�����}�ߟ{N�����t�??���;�Q�m��?���㞟J��*!����c9.���Ɯw�3�v�YC����;y�p�f��;Qj��t}�w���n�o֜���M�KB2��hza��M��Ÿ�\c^q�k5lg������5��}c=����<��>��ngz�/�Yu��W�zp޺:z��kz�޺���
�zh�o�5�0��ސ�M�l�NZ4z���7�u�ۉ���4���ۈ��ѱ�������GxNh�����N�G�߮}"�Mu�h���6�l�hy�'�������O���e�[7o>#-_��e�8ܛ���ۼ+ҵ�~zzu�:����o�y����T�v��ѽ1��ճ��7� ���������U����޸~v�m[+m�]���:ҫ8mKg��s��/�/��~oJ��!�r�27�K������>����q�a�_6E#��U86���^���mB7�n����|z�~'Zs/]��f��{��Һ����4nށ��[���M�������0M"
��� ��&�[�j���[���d�l0e�YPH�����B'%���,$����2�*�#m\Tf�%0,���JY�]X��d�B��IV�D��\�c��W�����>���}�<x�G�4>)��z{Ξ<��=��Ξx-�I��~_��z���ǎ���U����=�Q����=j��-�c����^��g�%�e���m�{'0ޛi����z�e���k-�x!w����:����ݱ���m��^4��O��>|kZm���M=����翡D���u|=z�==s�os����^�>������l���/#���l���>Ў���S�K���8>�g��-a���mW�Ϭ���ә�\���}��	�]��JF�����Q�l��+ύ��Z��/�-҉�{e�]��}���|���Y���v��ϴ{{�~k��^�<�lh��Y�O�m^���w�Ӟ�������}��Z��S��m�.ޱ��Eʖ��m�Ӟ��oz|õ
Ee){s�����'�ONr�n�����nK����}"�F[��q���}{w���_�,��~���A!���܎˂�>��r\yO�>E�u��'3��I�v� GG|������di������l��)0)pf^w�Z8��xZ]�N�v�d��P=�e��,�4����ReP�	=+��X�_�x��J � ��8]�f�q��	���L�.ʳ��੾kq����� Tm�CiH��EFb)�ե�c��S v@L�:Q���̸�	"�ʐL�AS�| �ܝ�EV��ł3F�(�>$���9Ȇ1��:QB�@?'2T��YvT�y���nO�<���۾�==o_�r�Z��o?t�6@�8��B����k�x'�_8�;}9���������e��F�g�l��������[��E7N �.*Pơd���H9P����qȇyex��T9�T��d���2DD#�"��J��<	���H�+$p�+�(>�ϜD�L`���E ��#��.�>; a!�vi"]GD-1�qg�=QӐ)H��$�H	xX��t��^ֿ�}T�X};����k���B��������}~�,�r2'e5(WNe'd���%�
$��I�CM$��4�őAI`��R�igOx��L1�yĎL
>CBM �T�Q.��
3̚z�2#�NH�EP�"9���I�96\��IU1�-���DЩ6�&�������@#���[7�Ԉb��'�aL���6[�%�DX�U!�'�b�')PSK�	C������e��ն:�P6�a�@��+ ��3b ��K�'4��- ����E�0���,4ې�+��Xd�1�(SK9�64�P|4��-�k*�a�Ms�J�Sf�����q�:;���(�s�[��T��m��dp��Z�à�iw'=��q (u�$9J�ZC�)���˂�IV�V��s�U4� m��p�!�0!�J�H���]�i���2	�55U%�n��:z��X�iP���љE���PW`�����N}��C?>����s���oN|[_Ͻ%��_R����>�ϩ��x}����{q�|�'H1������ߕ���딍~�o����҃����ĥ5<��)(>����f���"�5:N��m��	`���'��Q�# y��y�υ	Khڙ8���P�Y`bH���U��Tu�y�څT肒R���%Y�IQ"���d�eH��q�iZ�ʞ��� �l6���"O!�J�1��0B�g�e�ea��(�8��*���%���2Id�ڔ(�J�C����	�`����98 A�K���]�\ ���Tl4$������
!e��t���˥8�Bw ;�����G��V�p�EJ4��d��Y3�Y��3j��&7���>�o��gw�).�S_0�ٰ�W�?��	 ��2��d�ɵ� D�0 �1*-��5i�j֦ͬ���1P��D��(EB(��4*s��<1�����N�ÙAs+�ުQ�
�Y���?'2\��tr�v�O�;�`8˰:�1c�)�R��9h ���`Z(ޓ)�<Xv,v����������;���%:���^��Im��) �a*��i��V�Ć�!��j��j���[A�w�xYiFE�fɣ��!�Q�)�i��o�+L��\ �	�����g�qA�J��n	Y�,�r1	2�־��V�1ԅ� ���H��o.]'�3I�ԩ���4 }
lV��(����X�T��Xċ$��%q��׫D4GJ�^k;Qz�#IКq=�K�P����)A��t$Sh����E��DBB���r��RI����ʨ��*�7*�iMs�ȓ��_)��K�F�V�ݒqo<�0���E\[�Qz�&2�z��0p�(���V+T@LּIm ��г,AHѬ�K�S׾����@���-��7I)k4&��L
t�����C��_D�Ԏ��2UHzC�L(�H@��y�#gd�hҐܢsReK�q�,q�� +�$�-*B��e�)��^�Эw�$�CcN��<CVx̲s��!OJ(L�T��BC�,�oP�A�*s�M��}7+u3m�y��y��{�`q���(x�a!�9���
[&eb��GD5G��G��+ :
�3-.�^	`j��hÌH�u�@��ˁɃ���E�E�C�����\��A0�[09d�+j�j>#�R܈+yT�Z+����@2E�8M/d�="K��AB2.�*T�U�U�PX#<�.�-�b-�^
��H�"d9��\"����At���O y�� �c�����j�)�~�]�GV�kU��   yh2:���t��Ezj��CE�A&�3)� 
GP|���\��^Ɖ�c���\���8�8�&&��1�RA2���]'�SQ������H؆BLĨ)\͖FUi	ǃnx��B��{
�F����T%��C�A��YjjڑՔu���2Rc�V�,[&�u�0����@z�6R[9!Anډ�v[�C���"Æ��O :�5Y��2؀f#VB8�O2i�єF5�Ɵt�ch~��H��!ՓM`D��$�Vf6V��]u�@4!W*�F	60�*k�ig��!�$yA�P-�"[�ۊ3�B��뢸�@]R��*0��TBXm8xT�y[A��)�O�٩5%.9'\�pZ1�CT�LG����cM?\R�su;�ӕ
�3p"���"���&0���$�V92m��ah�	KO�'�U�7��e[#1UHB�	cf�Y���K4�DL1}!�#�C ,Az��"��+X�|����\/�����b�����
π���P��Ӣ:�,NF4Բ�J�m�Y+O�+Ld�0M�:�� edcOX%�9!"���\�uV�&C,�#��e+@�2�u�1XJotsf)401\!:eE�F�J�-���E�
��\������8\L�͠J[� ��":+Y+��B-@�D:d`4e�?m;$7`qL������5�=)\������Ud4Y��&W����!.�,�����8����`
\���$�?0�(��q���X���9g
���$�B��Q�,�2���S�ı"�9p��Џ&�`=E`�!���1�*��U�]�J�v#Mc JD���"�}���� ����7��ڦ��ֱ��Ս�� <��ú�kkK�iif��z��Z�숂�p�e��:f�.�-��9Z�X�I��I���ՒL�bA�0�v��A{�3�aB�h X#e�a�qt�
�Y�=5nۨj-ƈg'��aIrª���U\m�bbx�4�J�Q9�j�"�8:�s�R���Dd�Tg�ԉ'*9��A��*i%���G�㳌�`^X�sJ ��"�-MC���^��H1�!0�ȸ�\�<6G�30���j��Ұ.:�b�#�Cl ��+
�� ��ѵ�WfVU֜c5eq*�LL��AX��Q7�.-���;l��h(k�4M��'#-�B%�)!�P�
&��|t�8-���<4mH��KOb�.�n�Jp�b�p�D���.}Ro~V��̎�)����������J�T��4g���
�k�]�԰m�\��(�<#2��RD,(���6���^f�0����N���딦8�҉Qy��%���8�{pM��$�F�@ES���0���pg�.�����h�x�r�!E���E�H$���E�26ou�G\��XX�	C8.��Jp�-rL�_$�pw	�~�U�V�q{�ʰC9�j�eɺ�djS����@.-��~h�3.X��z%�<��*�,�TP�p���Ƈ78Ϝ�)��j�E�e H@�(�#q�>oV9L�&`�[RmxJ��A���&�$�b|��,�Lc�I����8k�'Ѐ��UK/"f��YHȊ(х�Mxe-a�<k��MefДbatD���Z���	��<�6�����
���se����R�Q�*8rnX	fWc��c�2MesC0'K�4�	a|���������e��p"��.�(�
����Pe*�E
��k�Zj�J��h�[i�)��Ţ���,[R�o&��U��\�k�\�.cE����QZ+nZ�m�5��mUU��lUT[j5���h�#E�F�*ܵr��+�6��F�h�[Ѵ4F���j$6���V6�e�:��ˈ�t�N���ɹ�F�t��1�\���o:�Y&0	k,�2�������K�1flk1��3j6��5T���B+����ADlT��"�-Eb����E{wRZ6�X��Mq*"�-p�Ii�l[	TTm��1Xڍ�X�6��F1F�#X؈�F�*ƱW7(��\ۘ��PQb-`���k%��j4fhرQi,Td�Jɢ�EET��H!"���?��_��x_��{kh����O������o�����?��~����(?c�>'��W�?��龼����,���#������_c������[�>���������.�彗o��>��p��|/����V��t<7���b�[ܟ��_�/�s����g��7;��{����V��������q��;�{k�m����xO���������-�������_�����l �L�ƣSHk�И��4�HL��4`l�Y(�!�1��ֳ6�61kXڨ��lTmEQ��QQb������`�X�ƋM5h��*M�������cI%bM�[jB1Qd&lZ,TZ�`��$�Vڪ(4[�V�ō���+F�S"ت+%��cj5�mX�Q�[X��ڱUV���EQj�l[j��mh��֋X����Jɴl�lF!4ADjI+L�Q�2Q2�La�)f�m4̘�d�D(&��X����������ƫ���-h�E[&�Uj6�E�mj-����6����ѵ�X��UX���[cmc[Xյ��F�E�j�6�lTZ��+Tm�X����mc-�c[X�TmFڋV6�Ƶ[�-�mm�+U���m��F�ZѶ���V�m�5�U��F�V�V��U�ZeE�@`��Tc�P��N+,
�,� �P|@@���^����=w����cQ����{M��|�����x����?g��|v����K��;�s�>���O��]�Wa��������}�_p�_��D��W��߯�_W�#���%�������}��;y�����>�����/����G��'�.�?����޿�g�=?�����O~���oO���������}w�G�_�'�������޽�~���~����#����������F��g������$ * ��� �*�]$Bb���
2@,$��J���H�0L�#$��ddA$&@���E2,f�2 ���!����Q$P�&�i�BHd��T�����$H�A ��RiCd$4�dB4Y��%#$X�"F�$e�BBd$d�Q�K)��e!HLɐfdQHR�3d��*!�bd���J4Xe�(�A��1`��D��S!%���#`�&$
,h� �04���L�F#2BRd$��`4��b1�aEL�2(�(`0@I`�f!�!"��JDA"fPFD$�IŒP@4��
!�� ����`&)��Q�)D��� ��� 2!"a��E"%��2h�1#!�R$%�(�2̈)��dQ�A		�f�2,`��bQ$�H"��2!���@4�Ɍ�bD ���2��P�!�&�F�eM
H��`��A2"�#Q�@&��D#�Ɋ-�H�bf2�2"ш���IA)
R��BFP
R��CD30�(R	�0FY�L�Č�d�Ѕ���I0E1�L��Ȑ�I��	1�Bd%�f(��Lh21D�d0��
f�2���X�?�@5pE� ] VAL`��g��|���Z�?�yϛ�e��G���w��|�/�}^��zo�gA�7���7�y����}�]��~s]�|o���?���<���7�����6Z�� RAT�Q1�A*
N�KAQ��N
?n*`]B�Z(�ـ エr� �_Z�Ƞ����*�"���-e1 
��DTm��bʉ�2�@-�"夠Q(��QU1Z��dj	PT$A[f�`AC6 ��d$�"9`w�)R$7�eห����s����_M��zӸ�}���]Ө�\�W����р�E�������k\����������������Y�?c��߇�=�?��_��>�����{���v/��~���}o��}����.V��=����O�컮�O�x�	��~<���޻O��)�=���
�c�����7�}����� ��i?�4_��澀>��{���O���e
��1����/�K�7��~��P���/�o��R@��R���0���EV��R���P��R�=;�La�%y\Jd� ����l阁�������O����pغ�ԀV(q��zvZG�7'�y�2�����':D��Kܸ�$O��+��.��N��B���0�7�H��[+ u�����W�v�jT��ȇ�2���0$8�7(&��u��4j�cbM���"����L���sO�^
J��.��6z�P=�B��},���<R�W5.��\��A�8�SkYM��-��2$�JXk ���/)~n��\���h�x�8.sc�vf�M!���<�p�yQ��_h�R�qe5`�t;p�&�LO��ۉ+��x<�F5F�w(��W�m
ז0Hɉ�+�M�,jf�u�u�NDr��1s�������㤪�� ���u�,G.CT�倜�Zd�b-1P@v!{��T9Qz�0U���Oщ.�Ұq�%1�i��J���q�S>HF�n��&J�%8_ͧ)W���G�@$s�k�������5FC�*"i��G�_^,�;���Z��uԠn8�*5N�,��4�%#),9�^���唂����Β��濌��SGm&8�D:����)�NT�U��9�=~"�Ը��Gf�[jab��6���~�H�1��K��B4yGQ���e�՝H��L�z%�};T�����3��c�Ȏ#��iG�� s.e�\I��X��W
�<��MJ�������G��9��O�pbΡp���/�aҥ ��\�;��dn�&�[':�����o	I£��_n���L2h[��q�2��4a���A�gF�t��l�vgEEͲ4��(8W�'*��Ύ��9j"���]2Nֹz>]a<Z���b@cb2<�0�Nj��
��+%�����[E�V:1 Am��.�>wM�(��58^R�;�0y�z�y�ƬZė�K���Hh�Gہ�W��X�@�ݩR��d�ѱѶ�ty!F�~�b���eͻ|Ϳz�e�aZ]���4'l[:Z��0�4�!��I�`��)�A��
�G���Z)��<���U�@�.��Y&�|$��1)�H�L���Y���㺕�1c��#|\"IX�����D$p���a]B�d���^�#h_T�@�eZ��TQ��%�d �]DI��k�\�u�/2�S-�D$�QjRIJ|3&M2x�<J|�L�g�8A�[���T�b�8bʤʌ��䡸�̫�E�n��!|� ��� �|�xa#���@|m�����Ism�j��{9�Z�W���og��8�کp�Q[Dd2@K�<�r�����Z9��u���+zmŅ#��r�T��,5*X�n����]�����b��3�̔�JJfg��II1�dɔ�Cȱo�� �U@�,�
���( �/B@@lQ�⠆�Qs"*�E��7�[�%��,?��}W��j��a8"G�5���!�Z��yBQxB#	Ƭ�_Ü�pWB-(4��4t��#PB�WQ���:��au6�C�.B�L)F��h	����]�}���ź#�-D*���.�P-.����\�W��6׋W��+�*�K@�E%�v�7SE.�䁒(C��.9t�k#t1K�2�d��(� 7A-1�1�.�%DZ�*��"8]��|���Ң8��H(�_[��ʋ� �#t/���Dr��Pp���(�+h%�LP�f"�U���DH����ˑ�Y��[-,��1AY&SYL0~ �\�����������������������������������xz ,���s���y���ޛ�=ao��7��G@@���D	QER�5�r��C �l�u����jv��RB!D�DPDR��{��ܮo� [ӭ @ ��P � ��( P  �     �    `�           3j�  � p  b�P�����kl-X�r0���+ڭE�j�������       4�;���P9 �@P(���� )��� ��0 �T  U��1\Z 
��M   �h��    Y9�\����    �Hh  $ Y�`   zL�姟 6   �����| `  ȳ��C�  ���                            �_4T)��  ��t�  8<�3���8g���x����
U
 ( ��
��U@H  )!T�P*�(�R���   
U��T P<ۡT  �  ʀ�d�ҏ�� (4��@�����(*�_>,�wpѾ���(�@�$ �$��̀ij�I�l;J�0�Ԡ������� �٠0����n��ERL�>�   J^W !� j�R�
UT��T�o����6�����v[`�� Р � O]�`%�*U�IU N� �   �    �� � >��m�2ES�    �  � 	�40Si��  2�=h%=�0 z`�L�&O@�	�0�� �4��=L������� �����&���C4����2=�hOHcMM ` �(M i��0� ɡ�LL5O��"�D�i���A�d ���=@  h4  � �     � �@      �I�IIQ5'�SO�=OHz��i�!������� ѣ@   �� i��F�  �(� �P4  RT�ɓ@i1�&��Й4���LQ��~�mɦ��O$��!��D��F'�ڙ2z����F��4x�i���z�H�F�4zL�*H� �   	�C&���4h h����& �C@4	��<M=L`FF  	�)��̝S�r�"�"e%iWK@bԎeds���[dFq�v?ztꢇ�J�s6�������o�>�c�)n<�?���k|\v��Ş���Ld<e޻X��V�E�/��ֱjE�&UŲa(1HY�D�%&G���|����?9�"���9}��{?JlmS�f)��1���?;�p��VU��m����)g��x�o���~o~q�o�6��5�����po��_/��{m9v��q��+���}�=?7���aG�7����7繈�vд�1L�Ϳ=?'��Tb}�S�n���s��3{�����}OS���65y'Zxa��Z�������)�Ns^��N�u,�v8��l��}�枣|Q�y���$�9 �!2{U8�s*r/�X�w\crύ�v@�}��vS�{gJ͉�:������5qa~������R�UU�����?ˈ��!D�h.�2MǗ�`"(�)pc�,�sǯ3g/t0h�N��{�����f�V3�՘@���g��qx�G��}�ݖ'$��i�x���@7	�K�	�q-�s�1u1��ֳ9����{ﰻ�t���^>��y��y�.}��qbr�R�*�"�i�sk��ݹr����� �Iqss�����v'��uH��eZb!:%l��&�QU��?w��'��������� /���������+D���~h�<�_�z�������:���8���q8��q��� ��C�����@��1��y��r���vH����ё�"}.��~Ȣ/�h�1&����Tud�)Jax�-��KUJ|�m\��|.Jh	�� � ��+K�I�n�ф�Q�Z�F0pdX�*��S��<ʜ=��#���JZʕC(����=��R{�<y�������vƖ�F���[�}]�2����2���f�(�����@��9�����V��M���F����$yy�w֚�i�\�[��Fk~�aw��$��5p�B�'/O'A|K�1Aa2�@1�|'֢�D���	SY�ϛ��x߄�P�l�������p��b�!�
(�DA ���0�aa.k���Z	����G������uϗ<wmF�K��LR��Tj��C�r� ���?�X��4TN��@�����څ�DN�kQ`MJB����7r�R��\Zञ�U�U��(��b�����|��>��> �;y���`Ï~3FQ� (��f(A�MQ����aa���f9������	�� L�nDa�����G����	
��z�0d�b��Q����Usb�]L�Y&��K�Ô(%�!2alO�jX��A�D&Bi"?�x��lDKd�ata�0�&K���[@���DSbb$���)���RjuO'#�?���ȝ�C��,)t�@�#c�
�Glݵ�\�8|?�ٸ:�,po��c7���6'���M�3p��\p��e�7�`����q=����u57�V߰�@ 
�SC(���1�G��OZU(Tq�i��3��C#o�탵g'z%9u�LH!1>I ��184�ڊ;��]LD[\�^�Q�4!���1�eM鄚�R�"p�(�AQ���T\�$J*�D��D�Jb�P �f��ʋ�(�NM̫2���:����(��B����=��u��z��j������O}�Ą��O����^��ځ?��S2�pDE����JC�j(Ѫ'U��۹��_o�@�U%U"��opj˨Ch��@8}=�?k�D@��z)TU�����:��� �����7���_{�dP�����z�_�)����x�B<vD�n��N�[�k�dKlR
"	��蹻��DŪ�,ld#(��D�j]�l�B+3䚶T$�%Ȏ�vlL���^\Ma�%��qEH(�L͕�̓E�1��*ؐfbR
a�>��cb�)
� e���~h��v��n̽�`<��2����>�Nj$�Q�81r�N�q�e7��x�y,p����M0<�K6�!s� 
bnJ���u�ٮP��~[V���q6����f��H�FdX R ��N�cEd͋P�z �*r �2"FAl��M��s�#<������M��gtF�A�T���4����Yrw؁/�Z���$��
?�V�����yy���������WC����r^A��8��p��ᷣ�83�q�ap��{��K��żo�ACw6�P2&AШ Y��@C7�n�M���ܟO��T�< ���~)��%�Q#�z���E�`v�`�
�������7�8� ��(�^{6��U@N���>�@R����_��w�G��o�m�b��y/��<o�g��d���E�s���ɒ���8�.H��[�@`�ꖿ�������h���?�7���z�Cۂ)@�D`�
L���r �DR�AY�16z�{=�t��9K��Н�Pe|�(�p�92��ˮo=kx� ��Ś�L�a�oџ�H~:�w�	�����=��$��e&�1G �)ċ����2���G�!�/jX�$Ce��Ј���q�?��>?x%�阁`⊼��>=�\P�$�Vߒ>H��r�����˺�N˂4F�/�TNJ�K]o"�SU��jM��N���!�7��n�r=s�����[���ѵᣅPP�H�aeN n7}�g|ߍ��͛��`����7m�f�׿�<��AX�&��)�d"���o�EkJPĭEBp�*�I��� �⑘�h���"�
���;V��r뷛ǷhP�̑.�ȣ���,2}�$�/��=����O�]���ׅۚ��PFN9�5m�nb��;9Ic��3�~g��3Q�y|Ǻz��L	�+������P��hiן|���Ӭe&h2)�!�p�1�T�kx�4]��R���[�eG�,^��*��-�qdw|�������+"���aR~���8�~��篁CCsEEEZ��Q�I��d��v2��}2���8m\dfy��3c��HA�k�lEH9�A�!��	��p
@!�,�Tj��htG72���:z�vA�Ƹ2�!��`��u0�Y#�A\��Ldd��Ab�g����6TS2��Jk��P0���+����,��df���#�O
vp4���0�0,(Ɔ_����G����ux����|6� ��wb-0�"JA)����QN���d��&��E��j��afh�����e�b�30g(�*,�%p���(��k!��A|��
�
zg9֢8���g�f�`t1�YR��7�F.U�vn+�A|U |�a��Sd��&q*�������ROЖ�^�+9�}����$<��@�`d��2�#�����̥�m�س�u��0���.�(r9PK]Y8-.*ɸ�A���NY�ŗ���a�����k�8�0M�*�l���F]�JO�Z��MT����cD��d��P�ej2�����2��b�� 1��C&x�L�������^3χy�4v���!�ڱ=���%,ٹx��2�\2n^xS�!)���v��JY~ɴ�߅l�see�,G1�[))�1%���0/�S�r��'f
��"��a��(@�&kCA�NWPkBJ�L�&�>�1�,��6#L%(��2���L�i3$�[�I�K�jM�mB{+�]d�Ft���K%���Q�:�s�6��l�&N�8CV��
qup��P��k��P/�%�<�+�\�ݟ����!�4'X���V+�>Na���Cy����)|�h󒬝�)L1�h.RT�WEHm8^f�k,3;�	�)���A n�A;(�%�H��39��71�6l����ڕ7l��Q���eei�NQ8��P���.����5�b.*��U�JT��ꍟ�k�����#CsG<�FR�TfJ�`�+�cbK���5<$���&��혌U�L^�3s���]�f"g#H�j�E���1�gG�^5׏�=�ۅ'���2�$X�x��=�'M%	�Y�#�([���V�eI�J��F̫&m�$���a3JF��Zh(��։%����I7gHZ��ԁ��P'=�e�?�W��ފ�&�e]�.>�}�rӀ}_3�h�2ل��P>N~{��ϓ}�!�w��T�Nn�g
��1Z��A����("��	�k�T�eh�N�HEQs��֭qS���ਵ(�,��h��ҍމ�"��������:��%��Tԡ!=>������>�s2qz~e~��9�	�a�>�Mr2��#�W�g���?S��5��Q6�
�?3�ř�"�r����ߏq�1�؏�D���R8���Tvʉ1ÕLuGU}G����!�~t���>�(d��v�Z�&Լ�Fa�:�	��FX�ֶ�e8��ԁ�����A�%�� ��H�`أL#
F�e�VV�b���j���+�_َ����	�w9گﾔ�� �f�f�����ϭQC<�rX%`�[\A�FǦe��Đ=�g��V��c�Go�3֑�<��z�����Z|�j�d"r����3�w�j��%�v�:ĆO�m�f ��8���D���͐���X�1�r�v��U��ϸ�k��QP��j��؊/��~T^ʱ�ܘY>�kD��,���0�#7�d8���$���wZ����u��ϳ�Ru��9��VK �SX%�o�N-U�:^�w߫[W!��k4��������������8$�TH� Ј|�	��JFЩ[�w�3=/�=������ҏ��JS0�3i��N���3cr3�}�s��^��{�8���{=e��
���'j�4��
�-[3-��dv0n�1��jޒ��uG�.�[gްYYZuɮ�Z��rm*��KM�{�4�zOU9΢�9��Bw9W���#[f��5�v3FقU��'�%���������Pη�g��j�R��!��ĩ
5-�ݧ��f��k,Fz,_�PT�1��'�����w~��9�����Zqn)0��֝�l���������Y��y�J�X� ��
��(D`O8R���%Q�V����p�Y�G�L,BE`�R�T�J 1ujծ_@8�R�:�1]��\���t����y(�rͧ�	�w8���*R&+�ļ�[��*���R'K���)�o;�H���Z�|��i����V	�a
�-I�>4��EC�`�!x�me��N������_���}M���1���붘�94���n�����mC���w���D{w�ߏV��Xy:��	8?�/Gx�(E�:�S#�B1h�5������
nm\0�1�'��lLˉh��>��7��Rb	C����Lǿ��i���__��w��Aȴ��l@��� ??�?M�iN�<���,�����_���C:�YX@,ꤎ��D5B�g�@���Ύ�8�24Y� ʉ
RD��o]~�����z����n$7߄#�����~������V��dz@ w^�� @f8�l'�>pd��&5�fǗ�:�%�b�� �B��P��P��K�	 �� 8�B�%���&�~�_�7��|�d�0~0� Ah�.��:00@�A �_(s*�������g���%��K4L��jR�����Q�!D�	�D�vBmڴ@�X�@�+��,�,�Y�1�9��G�����NG �"Ep@�`!�������I�t8}��%|If�"m�X�¼�E�GK��Mhق/�v��Њ�gg��J�|~o?�r/���Lg���Y�bC�ދ����!߷�-C	�-����� ~ं�1��_�n��r�k�P�[ce�}�V5w>#H��g�4b���[���1D�1bqP�0�%��,CbCY$3Q�kl�_�$�Ѕ��*X�HՂU��U�(B,	`�!����r�d�NQ�T[l�Zʖ�=bŇk�5���9F�,PQD@����++
Ņk[J,-�VX�J.���m�`j1����{ώ���c���8�i �l�kf��n�1� u�C�I�����j�z���Ԝ_O�Q�H��>�=���qi��!�7<�8C�{;���W�0`=(Q�}F�=�媵N�	L�Px��B~q{���>k���[�=���Cd�P�hܑw�{�o=���}����C��Ǣx1~��y}���{�j��{��<�;��=h_'y����5ߓ��d<�w�Bn���MA�ނ!?�-�{X_О�_������;�C��oa�J1��|'Ŝ�8�	�">j�ޅ�Bf����]���w����?�ھ�3�BI ��`������A<O=�P8��ԉ�䓁>|�F�N��<G�/�ݺ��H*���&���n�_U��x+���` o��{����ph�G~F �y/�����;��;@����D;	��W�Ll6���O��#���l!�2ժjӍu	R���C��?�}��X?��_�-� ���[�_�"�I���4�|Z�Ĳ&Ȃ���S����}i�}��"kNL���L��3W��ϛ��l�8���}������#Lz�,�C�?E*�!����jy~=F�S���f��*g(& �����I�4L�N3c�gn��z;k����u;����s���O��d�*>�� �L/a����>����s$����Dt(���pP����v������3���I��}~:�'L�@��A��lr�N=4X��Q~�^c�Uj��*����g����.l	R!�S����D�p��&C�j�Y�K7
B�B033#��Xw�E1JL�iS� �����{�Ȃ���T�	�h�g�U^�����S���Vm���J|���}�X�z(�P�����B���6���L`�(�A�Hgz���҈����|-��$����D"�RH��P�ߚ�y���r���>4Q�����F���/��E�R�ѣl
'��c�?��;�s6>Y�����y+��$������L�X� {,s�=�cZ��S��|}��~O������ u�L0m���$�}��ME�GT7l�,�фVH �d�91���&IA������55����2}&h� (��%�*�$W4T*"��!��+ ��dt]���产e�~�����'���N;���;<g:�;�h���rv����b�D��PNaAp,L,
BB���* ��)M�3���b��q\2#A�׼��H�����T��$�a�i3���+�Ι$libd]p���.ش���6�q8�ddi @��_"�rM����"ݜ�Ճ��!Y��=�%C��V٬R�r��#��3:�]97u&<��#��}�k5�2\�Jϐ����Y �+�)0�h�ٵʵ̴g���O�I��$3��'�� @�
�¢��<�
�g���Y�3������O�t�똩��_������%$$R�}���6R���A�$S/ŀ�jz�j�*kN}@�7�ȸ8���1���k��j+u@TNI���P�c�~�_��og�y�ߨ�a:N1��)Y-v��>���j�QD�b~W��o4�fK��M��)��J�`�g��vi�P�߯x�f����n�?s��~� �?A��m��Pk���d�0	T>�\�l���a>&���;:d�p{�p�7�QFB�ġ
�h&�x�2���׎" �ukZT���4�<�⇜D�+��aV����!�';,T���V�V-���1���
�_�����|����f%�D�쵂`�qP�I+3�]�(�W�٧eJH�³J�	�ZNm���VF����a�,���Z.��_�zp�W��3�k]wG�}\w�S�ڛ�}�{��5z�g�~bA5�I��社���&����{~eLe�e�?�'
�����J�$NJp����P�Vkb��bK��ݘ>߯��Q`�T�Χ�L�_����n�O��W����(��J��Fј�PL��&d?MB�����z�	<�pVsG��a	�Y0�SA��퓚HE�5���&豜�ԝag�Ft�)b�S��E�>�h����jy�Qq,&?Th#��f/�ֿ?$D~�����aIN_�JT�	.����i�>�s�j�Q2��?y�(�|����oF?������@���}<M��`�)\�KX_iU���Bx�:JbB�`�7��U�3��Q�^��Tޱ�g'�i:�2y)�4rk� 2�x�:,mlQ�BW�g��_&l�zG��A�������_��|L��FD"W�Q�Gu�g>L?�_�w����=[1����:_G�����G�n�;3��ߗ��F�;1���옚G{2	�Γ�~rz{��(�w����I����N+��e��b�bu��8�8�+�MO֌nuI4�H�J��V�L.�g����'VZ�8O�YYf��p�Yn���0+��W�8���{��p��wk&l�=�ͤ�K%.�x���г�HEi�ʱ��!�eX�J� i&VY�-J��Q&�U�5�N�5x])x30g�3�Mŭ:��s��Nбͨ�R�� ���ЫQ��=+�����o�]���^Ӟ�K6���#�1�W��ΆS�$�������-�)[�UN�ڋB���cE��
F�47�� �eh��6��l�06H8Đ=#Gut�e]H �dDQS;�����6��-I���E	T�1�B��8Y["�d�}�(�Aʤr͖�z"8F8�œ�����eɎj���c��Nm���D�	4��3DRIS	Mc�r^��4� Q0L%5CS-����>��w�7N�)�a��M��j�3#b����ic�ih��9i���J����ZZ	�J�����$�bF������H�"B!"
ZF& �bZ
J��fj��3e��1�lcM��6ͣ32����̌���ka�m3-��Ƅ�c)I#AQ#�ͫ��i���-<e�)�����(���S���3��s�"�R�T�,I�l-6m��6�T�TD��(iAPĀ&�g��=�:��.��U���
bJ4��cm�&Xƥ/=�5%�ǣݷ�����o^���x�z���T��V��H�P!� ���Eb��������c3X���)�Z�V�(Y!ajPԴ�ɅZYR�e&�
�°�i�mq��k��m#��[���9�_���r��4$0%Rn��35E
�A-T� �m���_�6�٬�����h��~*�Ѡ8���՞P���f�@���1�KCAKD�lV�[-R��� BDbV�j�2�ScZ�E�۠�������t�o��������u����h�Jc��jFF e�)iB��*�n65�-�ڛ,l3�[��k�|U#��!&�
�R��TQ@ٳq�1��XS*�5SI��Z�&-,&P3�CoO����Q�kv���~X"d̌fd"�T�B�-�� ��k�ZīJ�*"()!! ���<��d��u��_������uC0����V�"�m�l�W�-�ʯϱ!9��t�lq���g�hџ}�S_+,�Eb!(��b���8���nZ�b0��Wc����7)p�*��.;|̀`d�>&V�:B,֭V�����M�{.���7�C�vf�π�i�j�鸾��>~=K�t���������O��|��{/��9���N)޿?Ll@�9��z�\��^`�WG�3}ιG���/���3s���7��0W}ƥ�o}TM[�_��+�1��z9����4�t�{y7���/V!�K�y}x�E�4~��EO�u�tso�Y�o���C���5�+�s������/�[�Z�y��l����>oQA�[��s��?<L����̳���9�S��b�x��7E����=|����p�����1��q��m�:�y�u�k�<w�y"(�4�?��<Ձ��.l������'��'ē�I��G�������)̹�-w��̸%�8�	yږG�+щ�y��y.G/��wiS�%�y/?Ǒ�wq;���u\wV~]�.����݋ē��^�O-�O�x�
/'����?#ӌ�Y�^�����v�9�T���]c�&+6����Xn��uSL�x��ͷ�}��v}y񶻐������0"9�%Y^c}�i���<�������6����^���@o�kʌE 9�����]�r�Gx���LBzIT��Kc�W1~X������-��[�߈��pz���.Y~����y�8�B��\(�wq��9K��O�����9�a��U֙�u�{��H�]Ψ+��~#̧�s_��ߓ����|&��m�\�9���HG�鸗�1�#�p�W���s����:%<�H���FO9��~���Vn��C�l�����q\we�x��z7�񜌾BO'����/T;�7K���d-����K�܇o����|���,���;�p�|G]s��%�j����_�Ӌ�����'���9'�.쾇��1���-�w¤���y���?X<砻�rD��I~�?������<�=�wK�~\Vp�v�T�Y��87:*:@��v�֮����`�9�!$r��K�k��������/a������){����8n{�����D�.I����D>��iw���j���U�a4c,�CWv�XƷ��_��~�*��B_��Ȳ}�20@�!  RR  "�L>��5*jWg��\�yD"t"  '�<��ß-KPs�76H�[1�;�72��� �`�J3\ϝ����9�R)�]�������h���@�����a|�!��J�@��A0C� EKg�D��?��	�D(DBu�t�k_��/O�q��Ԇ������j �s�M7����
I���УiW����z�) D@q 
"3��l����']1���d�DV
{��S��zEB{�鑐 D ExKu�7^�#ˇ�[Br�é��o/�Ӿޜ>�@���}8i��$�l�C G�<���;Dx�I�_d^7m�߿y߿Q�0@��  `��E�{|�S������\�r !�@�DDC�Z���v�-����0�5��������cEh{������ˡ?O:��1������Kx�K����0��~Ǟ~�
v�cs�� :@H������>�O��?�ޞ5��3�t��M]��2��ߔ�iلs3��W0@ 2 ^>�.��{�� E���x�e�u���3�0�c�t'�OƔ�2l;ŷ�p+�]�wt���K����|ϷOr" �@ ]�T��$@l@�q��ڃLsl2(�jHP���>`�3�0 6�K���<���o�]�� ��.���g�u���_J����,�_��7�^��<~�y��RQ��o�(�><���c�zR3�/���@�@ B��}k�,�2��~~� �?��C��Z����v-</�wc�d�N��x����Nq}ۋc�13����$  �4�i��Ͷ�ϳ$}}�z�h8�Ѹ���r�1��}�Xി���Qϟ���zˡ�yx�<�)B��D�,q�k��8�.������w�����;&�}ۧ�}cwe���Cײ7,�^������ �K�j�����<=����� �J���;q�.pf��}Y��� ޱ�6�r����,DI)�oȵ�p�9s��{���D� @W�]s���8�:Y��� zq?��������O~�����ۇ� 7ʳa\�v$��x�Y��\\`t���#	X���)�U������O^yW�� �Ig��V$e� �*X�'K��Z&� ��hLlC�p`��G\|�F��y�u���?PD[#1� @<������|���}��I�����~��6��� Ld>g�}�DJ���Dd@ [�����ǎn�}����Xʼ��� ݇O�_mV�c����gŒ�t�Z�<辰���
QG��7����_r��b�Id�_����y�iQl�"�6QCE�����!F���{Ȋ��Iű0%#����ͭt�%�E	�uJ/��:E[��zq"H�u���m�}8@4%�l��O�}�~��z��z4(��3
M���,�2�q��1m�B��"=R(�h ��Z�� ����\o��k5HI�.U��<@���������)�R� �A�k9����� �8Qᒦ�/���B"�X	@ [��ޗs�׊Db1�������C�Ek�E~��A�t�������Ԉ�",��-�w�> SښCG�ojl9f�/�@�����C����(+�윟�'�֝�C�{�����}�&G�|_�̀?�ܬ߇m�{Lq Dx�ƾ�n��+����-��!ޕ���s��+d��ϗǤe�&�t����D_h������ϧ`A� BDDE����q�Ӓq��d8�ff`�u���?��B>)|}01��NǷ����0C�ݺ�5�������D��@6�M�*�>��Q���vV��
�M�����@��R*��ؾ&� }|�g�O#�}~����]<�� YWN�3}��e3��[���7Yy^��i��ݟ>���pf�ye�k��r{v���D@�>��b������<|��ɶ�Q<��r�Ӥ6�n"g*�M"�x_���x����7mL@F��l�h�)m#�A��D
��t�4_/O?2""!��)jj��?ͺJ������n�EFf�D\��(+�(d<c�2�.�T�u�u�j)*�ŬĚr�� @��|����A�UO:�	/S���~#	Z�?Gc�$Q�="M�.���0M�D��^a5�4��q�X��J*�@z @2"B���M}�����e���>�e��r֚�'a���ۈ � s���� Ȧ�W���Ӿc����/��P��<�Hմ_���""'󈡱�6����	���"�@�22/N���GӨ�,��ƈz�����RȈ��<��>�A  ��!���Ll���]�=�9��r��T���r�oj|�?��*>����cg p`�"��Za��=�ǟ�U�d���&��k4���z�n���Mv�A}x�Ν������3������	�h���e�j�����}�v���>�E�9 ��f�T\�Z�P���3�:V���?N� @�g�ך��$�yqm2�3�"��գ��ra9>͚m�,)��A$�q:h�@n��p���_�}~;�� 72 @�~u�˲C�N����i��Mሇ�M�zm��h��au�8`oxv�}�~���?JW�-93���	I���;|��s��}���<H� h@� D4����{�c�5�DM��<�yD'�E �r���Z�Q����F��xsK��Q�2��������������|AY u<�wWߖ];\�Q�^���ƴ���%F%�%x�����@�b��6���q_q�C]���]��4�O!l�{ @�C�J�[�|k/+����%�mU�� �����9'�럣����d?��,s��v>���e��A`Qx{�����x���z]4�-�e����yv�E��CHM����PE��D6L�d
I-��}V�Vd<� 0@ ]|��TT�H��+��-i�8_��s���������2�e�q�DZ�N��;c��עp  X����t��|�Hs}�M_�Ñw�k.9g��x��p�/[�7��z�Yq�4����(Ho�""" �I!�d�9�z�ٺ)���*��w`�i PSD,  �����R%p���i�����o�2 s �� g�����i��xJC��T�.��R ���VU�`�_���z��B�>M�z�>V�R?]� �e}�W�\�yg��+A���ǹ�!��0�߁=�����~�?˖D8ۏ	}��;!P@�x�A�{�͑�ٗ�_�>>~<�?���N�����ǋ�C�}]�qp|S>�~���ic����۴~��9MR>&��5��B%@hdD,�D�>ir�.�:�Edy�_�u��%������{��/^}��8 �i�/��.��˾���B܈ 
F!��W&S�O,�r3��ʣ���r͘HG��KD����Bg�e��{� w�%T���	������t��,g�oh��#,�3�C� u d P��!�+�-@ M��(yk	®$�޷;S�����s�,�8T��}z�֯���Ёs"  �0D@����V�e���'HC�ק��V�c)�v�R���=E3�xf�A�@�@h��.��}O��K-n��ӌ!}��y��������yG�]>6H���7W��JZW���Ad�=��62  .`!����Amկ�$.1�����¼����.����Yl>�>��B��f�>|��=�n��Jt߀l��Ǵ��" �Kj(p�Hӳ�ڰc9�ENH>w�M#e�T��߿�1V������3���~�!�R�T�^ù���'���5����/NV�6ɺ���l,�ʷ �{�Cf�5tL�����;N���=���dDD��y���-py}zo��  e��_W׿�?�x K�:F������'�����znC<�䁵Ƽ��Ŋ��.����.���M{�,���Ғ���H*2�������.F �3<�Nu^ǯ��4c�܀ .������#hp�w��-Zrm19<�,�y.� �|�*O�G�}}��S8x|X���,�N7H��|<��6�M>w�c�#�Td����l�iB8Ǉ�! ]�t��˱����� �<���o��ۊ��-n"��G��F+����t�!�:oj�QBP�d�.� M��ׄ�g�=y����r�@R�S��'lrO����b��տ�M>}|`��g�/3>|�s }��\鶓��@�_�"�#�?Mu��!�(wu�����������\� @ i��闯Nܻs��x�c�d�w���UuIR\�+���m������_�ݙ���j�>�\Զ��[�ػ;Єh.M�0��mǦ=�J����W�#$������'���ڂ�J	�v�e���s�ؼ�i��ZR�~���^�K�\���}ei�o�ހ�>JՅ>��?>8ڡZ�M8�u>�o�Y�����~�A����^�W��Ƀ�u�rh�t���}�����P�c#��wwn�NM=����Y#l�-,����|��ZP��z֖mh��Yy9����5�ƯR��L�̩����3�bzZ#.�7%s֦l�(�������ۏc��m[��;v�^ي��������v�[-���k��O`��v�9�o�Ң#%�n={N����Q9����Z��Yk�'��q�ˮ�Z&��iu�uQ���6�k�Q�jT_%�+QG�A�bεV������z���y={�t����e�s�Q}ج�T���U�P�Mram�]����u�2]a�b�M�OY�o'����uG:�Q�����y�Tg�;!����Xmg6����.��s�* �*R��͏&����ErZ�E�.��l#[��>���	�^�F/�ȋ����*mA�����䵫������o�w�p���怹G��J�\�kR��ׄN;V��ckz�[<��K�Ǿ������ݺ�5|�8�Lf��[vq}f7i�TJ��Nxy���ֶ�Ƽ³�|���G��_>��ORy��}��<�7�o{N����맟�K�8��v�V�6��ze��K�u�4��
1����׏_3<�n�uy�����cf�����W��5���S�:�Ϝ���g�y_����j��w�o��7%�i�X���^�d�;�P�+��!g�J�-K�����֊�Mv���Z���T�u���sv���lg��;wQz��JͶ� |�g>;d�/�3_!�o[]u�C?&N��6��m���L�H���Xd������(�4˜�T�����Ƨ�TomK�}y��M�.�v�eG���V��/v6��[i���m�z޳�ϻnݎr���l=�]>�/�p��V�s��>�{W	�;��R���-�SQ���v�gnyS�O'3>�U��˾�.�͇~��z�&��%�GQK�J��'�z�$�����QZ�By ,$ ���w�?3�} ���[�ށ 	�H �)	X@X@��<>������L���W�������i��/Y�~{�\d��+�1��ر���]ڕ�;�өm�A=�"&�����;v3�?B�%��[ƶv�[��b�m96�����Zu�������T��Ҧ�U5��7��O&_0�j2��nK+�T�<=��e��mg��j.>j(�-�ZE����װ�_5�ۅE�L���%3�S"���C8i��g����q�f�����o&7�Ff��?f���w�(,}��N�o�V�Z[�듭�<�����o}=��]��9(��R��W�6���iiA�O�ǀ�:g�~{�d��U<�v����f���{Oz������F�����M~��ƽ��"��휜�u�Ue��;�\>����5}�mDo�˶�݇�䩫T�64iQS{�)��z��%�Z-'��-�[O�1H����qc�C���DY�U_|mO#}����޷��D��څ�u�n���Ɲo��{���"H2	�j�ɩ�fM6Xc���յ1��d��k�,�j�XY��1251�E�&,���ֆ���#�a�e�1\m�#2�jшښ�e�Vj2����#R��fi��թe�Sfe����YM[R`ZM��3E���+ZA@��!IH�.lZ0����ڽ�_�Q5���m��k�V�E3�BוÑ�N��ȥJ���{�������|R�+g�Խi���r}v7��䮣E���'2�~;�ss��]+a�MG�Z�=�m[^�����������8�{{�J�o�Y����^;q�����X�d�h��M2"2�q��^��]N���k����z�{�΅�֞��Zԩ�o�������׾�����=����m�vl���{��N����w��=�-h�>}{��
%��>fc�W���L�-��S�=�ʫ/4>$o�Q�meHߛ�Z���Qg����_���}k]�C����Yy��ٺ��'Zʔ����+���s�Q���L��c�+�J�Wz��MF���(aU��=NGu�ڕ3x@{m����-o��Lj��~�?>�ߐ��J��Է�mz��y%����;�Z��;���n���޶K[[�ٲ���J�k��YK�5����+�*樣�;��~�6��{ (��ڏf�+Z����R�W�jV3���GZ�䢇��0�˶iV�b�䮴��{��B���h���9�[nTQol�7�m�S���E�j�R��v���ݶ��T��=�2�k
�k[W6��j+��3��Fq�o��Q5���-�^ݽ��ҭj�*,eB��,ػ��>��jz�v�~��z{��My�����E�͢�G�Om��=�oiE������Z_WrS%:숛�a�Q�[E�B�ʧ�{�ٍ�+U���24����Sk���ѧ���Ŷ=��sȪ�S�=�^M^����8��e���4H')Z���38_Z*Z_����\���B����l�5��M�̕��o��M��*E������Wޤ�V����n��5�̋F--��gOjk�Y�U�o�ϯ�N"��aG��[��i绗K�|t��)�^o�(kw<����,���m�A��A-��W���T�cl�J)JV���}������O�W1��)���]<��uV��
a6j��7}%�֧޿wn�եJ�&��Ok:5��l�\����n�`�w�}����i��r׷�䴹�$c���J��!�z�%Z���m�J8{�TY����X�Qo�L]h��ͭ�mUmR�4*|}y��_�sW-)�R������sS[���g5^��T<ѯ�����Z�&V�m�(U�=�wek�s9�>ן��u뛦����8EUR���R�Ľ�u�v��'}����Z�>����τU岖�b�T5����GZ��Q�-�S�L�%O�?qϽ�Wݵ�g�_=�s�sڼ�;6�DEOY~�����KO����b���z�Q�l�5�T_3�}�p��7!�s;��+Տ��z�o\�K�;��sL����-���j�;��l҆ J���>O�*�}n�s��S���&�jjW%��KCb�\�}���͚7�:��+�Yԧ[�(��E����69��Ϸ�n����_��/!����R������u�mcQ�K�WSki�[�SZڜ���k%��K���c&�ҙ�����U*.ˌ�f��]|כ�ϭ|֨�6��1�-�{�d���E�G�o%Z)l��
0�j�_q����V�}�wk�K��}��[��5�|Ӌ;?]��R�1]=Lm�E��"V;���m���)r/^�]ܹ(ev�Bk��=אo�����>�5�5��/ֹ�Ylgu�Ӿ�������5sT����όm0��ݶ�J���m�E�SZgoq���{���:��*���V�W���!��*��\`���Q<	����4�US�R�0�Î�\(��)*md�l3'�ͤyL l���X�fD�)HIbG� ��	q&1��	@���=�Z�TDZ�X�TE�A6Ԩ#*�-ab�`���?��`TUb�QAA	��������[��������G���8�� �<��[�;�<�f��GuVfw����,�u���k��cc�v����λ�ɗ��0r���Om�l��EX�A^2��~����P��9|�r��~߁@��$H�*��%\.3I��c��KEC�t�q����&2��b#,�V%U��xݞ����p���8�{����� ��f���*��� ��^�c�9��%�9�kF��q(�}\`L���)�i�ە�;J ;C��"��ҕO�)�`�������Ӱ�M�.�_=��}�^�eb�~Ƣh��d�R�	ʄ�0�)���%7Ly���Io
�"H��*ւ2!�\L�ۮ�h�,AF��18ɘ#�x�Fv�˃
�{{�.E<^^��.�"��ύ��1�2Ȭ�ő�3j�+a�����F'Z��5����qՈ�5���14l������E�D�;�aL��Cxr��"�L�)�R�Ή�ǖ��"�m�~:��l�А�/D��Kωjd@���=c�^��=�K�Cِ)΄6���Ҧl�гe��7�Q�E<�0�اT���=mF�#~��l�d��J]�Q{ �%(�)�P��R$Vcxk��ß���0����Lx��=-Z1;z��GQ ��(���;+���+A��\�(9��A$jD�xtFKnf��4x����:"b����9�|rh��bh�Y�x`H�c��	Zn+}��ZW���۳Ca3�E�
�+c-e��G��7�{h�O�wafE� ����V'�2���Qթ�A�!\%�8�OZ,M� Q��{�f�|�`��fpq�})�G*�o��8imrFU�4���D瀘$�c���.0�1֪X��j�	����)""�(�bR�jj���"&(��(���	�a�����*�)�����j"%���"Bf�b�����*H��"����" �)&Hh��I!������b�*����*��& ���������F����8���0��!�\�B ���"��$?����+��@�_��`�Q5A��h�`��kZ(���Q*X�[Q�X��+"6�V�[J"D
��E"�EU"����Eb�KV1m�D���m�T�QDQaZ�X�Qd�*҈�`T�j*4l�`�P��F
���bQ�U��(Pb1��.k���'�u�2���y�O���v{����ی�<�)"�d�~�g�������(e顿R�)�~�r�O�c�����؉�L8?���)�����jH���$!;�w�`���0ia�C�����hǾ&.W�XT2�t�Ɓ*]�)`,�Bf�j˜29ofSY�z�G���+.�pyn].��CS	p�M��7E�0@�fr���k0��.0F�#�tYBBG1���;")��f�;0w(����A���ܽ$5�[+ׁ`=�n��ʹb�^{Ԫ�!n��^�IA��Dω��1�v��+L��Q60�-"�(T��9�\�j�lx�εe��8LM�s�	XY췇N�4���Q�1���OO�v���Z�7_[:ȍ��K���ܶ��KM��]�1���@��/��!t"B*� 놃֡�Zt�I@�E�5�,�
�w*/���ʇ��30���+�RN�(��zњ$g;3v��+��s߲8��Y�ʚ�7r���2	<�W�luMv:vʩ6j���:�h��~4�!lQ��SH���8t�#R��rH�DXc��U�1$;�X��c#b��ڗ���D�H<���P���Nl#+�
�14kߎ�N��1	���7���a%!ҳ0i�5����K�\'a�pl�jj1w�S��i��<�G+w6Yq<l=�<4Y��3�I4�<%������Y�ь��ՙG �ڎ��,E�I
h� 㚖�qX�o)�6m��R��F��z�i*��5&��3��F�A�m�P�����e�/�ނ�V�
��{H��3 X�*Y�N-��ƕh
��7�!I���N�7^�#)�)���c�6����5��z�Q�S�^������m��bŉ.����6#���R�ŕEL�T��"��4�d` .�t푏1y�
�P�G�5�(JLמ*\%��m9[3[g$t�.�/�;��,�2��Ʉ1�yxp�Y�R��f��I�6�o��d:$3� � Q'�ձC^l������}�����*�d*�U�j�4��C�ʱTD�4A!M�S��SRQ���IP�PECKKV6[)�2qy:�-��� �1%�\cNA}jx���+UU��H��,�D��H؍V����-���X���
�E�5��ր��+R�c�0.��W�z��G<N����j���ʣ+�E�P˭�F�PK�.�����UrUEUE�b�D���$��֋\�P��Df1L�m�ŵm[V���E�Ҩ��meh��J�i��.ZR�5֊E]hT��GP�3X"T*�U�ژj���k������i�X�(��A���'�� h���CEMDPUQ$-D!E4ST5UADTSLQ�34$QEQES@���D�ci&jڧ�T�U�/��U8g���x��4��w�u����ap��N6j�TҀ����
�0D�Im2�ь��4��Z�,�A�F�$��=�BBf�s#�����B�%T��)�)(R
I�v��F�P����ZU��E� L0G�4�6~���U�l�����6 H��,��-�gv��*l��M�f�5�4�������4���*�Ύ�9\��$Թ����s��&d4LQ���}+�����O��;�itv#��W�\qr�^N��r)�}�9Ӻ2#��lG-��bR��ؒ�V-�3B���d���DrD�CWOI0*3��ˉVe(+k�4�,T4�P�����r��y�+��ʎg�j%Ip�:2�7�����'~%�L'~8�E�X0
���@�`���8yKI.l�i�q$DL��ܜ)�Z�0�8�n#����	+vS�2����b�J�@O����*ZR�~ؒ>o�obqo����BiI�:�y0H1-4�6S���p�:�ͪ�"��)�:��Z�+53ת����%̜��j���ڵ��(<(E�N}��:�x򜙌�i�;�1IJ��M��v��O~R�)#Z�@��K�
�\��q(%!3*~�I$�u�B�4��#)6l1�i�n�ҝ3��TG}hxJ����R�fTy����K��z4;�8�\����;M��-�����ғ0ЄCIHD�JUH�U\E�Q�%emQ���q�x��y'�p5Q�;:�7"P���G����g�ϛQ4�V�3p>�����|/�?���v�v����k�f��M��;�3[M�
����޸12�  �?��O����|��C_+���G���[��� �����?f��*_v��zYjP� ��;m   ��w������>�1~���~Ӱ��l����~�Ӧ��[��W�vO�ز���i��������w�-$��D3e�7]�(d����#� *��w�Q�9/M����z�o�z�����;=��˽�;��ѲϜ�#�T���)��䃁#��~��}���?rW� ����k,��0}�+���b�U�!���?Pa�^H�kg��^��z�q��e�#�CS%O�������=��5�ؗ���ۇ  ��3`~����=!�@�pYc)�J=w�����r�^���T����;��Ka�`%i(RIv����E6�.f�%3�623X]���ɋ��O��i�=wLj jʊI0@��z��e��k_�v���s瘤�C�P�_z��Z��KR�&-IG9��l�uQ4@ۯ]�MP���}������fϱ��,�6>j�ϰ��9�m��:1m�#���s?�Kˋ��� �g��@Ƽ���6�Rdfze��O��g�n7}Q@u��kv���l5�����f��|m2����d�O��p��-[@ւ �� 	>!��/O�#�Ɵ����#�S���f̘�r�'I�n�-c����(Ca��ǉ�J
h%8m�2�6�%<!�[=����h
�"�֜Ek@��B��]�S�P�)*�I ��$#ґ`�H��X0��@�\Æ"a��hr��t4���͐�����m��h�l��"�b%��ZQ�Y%�i���U��UZk�L�W�Ì4��#b�
�9��<JPl�b�e����=������'�f(D�c1�ِ��Ê:�l�7� ÒTEdF*��Bd�J�� �	+ �I ���w�DPam�Q���66@�JڛM�6bF&���&(H�ĊdVE"k�@X	�XD�����¨b��J%'��&H)�R>�C$2��mh];<}��x�[M�X��)	"FT����~��C6��l�6���q���y��H 1d�� ��O݀\�@�(6����-��PP��Hs ���� BPE��le~d�!����Qjr�i��nY�lh�RM%(�H�TL��g�y�0�"����رm�F��q�r��TY�e�c$ Ԕ�ج� d�̩
0B��E"�	U'� I,�F	��3"C���y��f�C+ejf���EN�M*�i)%����Ƹ3�qq�հ.��N!�s�W��6ɰh��d-�M�N-\�i�+,�ۖQ!>cKZKa�؍�mV�	|mhԳ#b�C�f	4�T��S`��UM�mRl�[
�eF3#Cfƭ�=T|�S��HT����:��$���T����?����b���c̞����H|��b�';��UmU6�����F�Pڭ���[�ت�j#b�$�X�Z�U$?������+b���3@l6$�cNY�b�yE)i�bi6VjSb�iT��I��"�YUƐ穵n��b�C���_'��d3�Y9$ ��ZR�aLn8�va�C�-b��&}��Є�����侺�jZ�T��\�3�c���F[�;�kid�u�wvpM6[@:�p��B�p`7�g{�g���.����^��-�fw�t��}��?>U1e�~�n�+��gw��Z�=N�L���PZZ6�����_p���'�x�������O�ն�/w�y���m���ž�ox�kS��~�U�''�<�C�ۮw��?(������m-(j�^���(}�.(������ξ�h��y=䳪Պ.gɓ!ÕU�����Z�]��S
&oWT1�����=����|�2����5�X������bɨUm�S��������j9G�;`�Uu���Um�zؼY����O�q�_���6h���>��KlG��/]�ڏ���5���ʉV�Q����Y���j�}z<�����u�yh�o7��Z�:�!ʝy�ԿR��޾gu�[�v�~�1�wl=o�wK{�yὰn�4c�L���U�����C���Z���X�w7{p���=��~����7ws�>�c���c���֙��{4�S���}]E�Ѷ&�1��ƷU�R��n��k��ɵ�����ǵ.��*���x����7�O[����]�{��潯v�Lf��<�q�2L�gf�JQ�]�/�j7͟{�U�R�m}��J�>=L��=б�ݮ:��v���A>����1��֨�&�����l[m�{�����6ɻ���\�l��\e�l=6��wޫZ9�v��}׭�c�y���-/V�Sam�����>la֑o��M����G��J�l����c�����l�b�j���o��Cݼ�n��)ڮ�:w��\z������ë�lY��|���Km�L��|�&Ub�o��}o�:���%)D�����Dz�6�Qc���7nxO���J�e��Z��eQ�ڣm7�2d�z�T�3�v{y�9����i�;��{W�����m|�Q���<�>�"��QK[�e�������4YM�O����׍w�)�V�X'R���oqrf�{`�gf�j[^q���ֵ�,�sb'�Y��o�f��J�Z1]+m<߯�Ӑ�����(�}omD�~��m�~_sRVE�U5eJ�[W1nm��2��S=oKc������a�r��[�w�f��e�����Q���h֭��3Z���K������}��.q��۱�h�uw�;u�%}�¿}}�D뜕�&jT_9Z޾|�����
@ O����� 3�=�@�����d&�e]Y*���K��G�J�됕	<��3!� T�䕒a%IU��VT	��q�ݚ�jGV��ta
�y�V )� ^��L���|��Y�,r���R:i��9�5c�e�e�6X͏���zo��4��F�W��>��z�wߴb���w��ƣ��<hŭ�̻W��bn�ز2�Y Aa��@�w��ߗ�>ݻ�vo�3"�.���<��(�?�uSj҉IU3ƙ�k��~����^g�j�\����p��ϻ�d&k41D�!`b}8e&�T&�7� {vN�wv�|�?������?��k&l��fͩ�Z�5�(�7�Q�����'�����TU>���
��*Dz���8�x�&���"��+6�
�/���p��5*j��jl6�.�+C�M
B.'4���,�Pd))�"��'���M!J1ACIH�ADIKIE4��QQQH�EZi"K4ZT��O@�
�@m���"�M5b�4F"Qkm�b%�ڱm
"ZQ��)�qb�Lq��}Q`S���χ��!�^�<ɧ}-5
D�Vt'ql�2��u����U4u�I�����O�����{���k�5�k���A�������K��=�,."�QY����Z��v��s5|�1k������dE��x�C_w�i���E$3]�ט�[}��dy�e��Ҡ��C��\�YC}�����	0�␒��ܐ�2�S����m�bъ�~���]LY��}w�C�V��a�]�e�W�i�g4|���r��>G(h�|?!��W�n�m�6w]��D&�cz�J���s�7��ޠ>��<fק��g���/���h�_{���C�x�����xޙS��Ow����]6����@6������}�C�z� x!�*�������ê6v'��|��]��n�~�����>������9���:�Q�{����Yj qc�O�վ�0|N3���</yD|����Wa��֟���<~��~0=��ы��K������oY������[�������d��HkJk�E�sz��) z�9��K�g�e������f�yx��@	FO���'�d_���{�B �d"7�����'��\����!h��|���c��h��$��1)
��Q��j��!���`y�r!3N��q�q�ӫ���>:ǔg�2>�1�A'W������!����ܸp�V�/ϯΰ��s��o/�e�)"i�>�����R����ۻ�{p�A��JǄ����g�M*�:r�//�������0�ɡ���|��	��lW�O���u�L|�XF>o�W�5��������	z�>g3qQ^�\TD2n�)彥����3��O�}����q��))�Lx���rS����Mt��'O�j�rrF40F9�	 ��*M(c
 !C4�	B����a���H
�q��-w��Y���)�{���s��idߊ�
�x��t�Q���o4r��cC��n�g8����iO��}bʺTD��t�a�n9�����3z���Gg��c4ͥ��|e��<i���z����I�	2�n[�0ƶ��o�f�!(���y���a�]��z�e��}����W��3k���(Ҹ^G,,�ZZ��6�|���M�e84	 v�XZ h΀�iq�$��T�jr:0[D�`n�u䱲��GN�@w��6r�	3>�N�f�/�w7dr֙�&���8�e{0������[eO�}oX��~5�H��虹���X��f!�\���M�d8�Ù$y��������uJwSO����/<���/�Ͻ�ׯ�1��i�δ��ss��ɸ�^<��_O�ɷ��,S9b3֭58i��{�ק�f�鮬>~�����ϣ��ڑjk���@��"ިȞ��L�b���^��ib��#\�苽uޥ��F��Ä�̺>���(Jz(��ԋ���'��9���� ����\�����e�
�jl�jҶ�e-�mEl�lR،ʫ`�b�6M��6S��mJ[Pڤ�M�%3-�,�Ʃ(*i�&����J
���������� �������$F(�)��X�!*	(�(H�Zf��RU(����&��me�l�b�Z�c�$�*#jD��![A6��db�PM����d[ImTm)���RF�I���D�!�2b��s_Q�,�&`�a�i�-V�m��ښU�Z��Y����U1���H��ш@���/KHH��m���W0�`ˏ-��rϥDj�\�G8;�:
�8�!BJ����*Iai
�`��b������+�x�.0s:n)@���WM�J2I�]EA@X������
�W��I�eWA
%;h�3�� �K����J�
Q
(��B�3�R穴FҺ�Qӣ�)`��AI�������IF��X��A-��Z�QY�=h��T^n����Y?$��2:�m!'�!<�O���L2r�*J�"Ո�YR�Es*3*V�E�mAPQ��� �J1UES����$� C�%@�"�k!��(Q�m�K
Ϛ�XTZ��YR�iE����b"��"
Vj��=աו�z����2*��AAf��dUD�QEJʡ�p�D�J"�2͛!��(�(|��͹��c��l7�9z=mˣ�~O�g�\o��/����5�����=>���-�s�oJ�U��O�����OIȢ�%�-acu	[�CR�����Q���j��*�R��a	@����EH� � !ȃ���g�%^6�a���&�B'�4���g����o��_h���]��yr%�C�E'5�#���9��#���Kh !���(��O�d4�EW�g�=f�AE�,��%�
�������A�� XT*/�(����8eA�PF"j��U����bVT���@s��$0�2��F!�7��u����魸��W����v����X}�sT�Ư��!���e|A�[2����9���x��ƦZ}�Mn�vM�/vRUt*�|W��G���7�I&��M�{������Kc4���3l0�t1X�h0�JiB����`���\�I�5�	�S,�H��eWT�l}*#B�ѹ�����<fݣ�''.F��	�U�q7|wp�V���&��+�x�&��d/�P���	Y�ޫ�@�@JU͎�6˵Mg�t�D�	>|n���Y��j��l`�P2F�1�5�M�u
V�L�d�W�jJ�wek�ݍk��Z�b݉ۙ�b�kݚ��P�d�n���̸��ʲ��@�5���طd�]q���t^Ц���}m����ld-�a��N���Ҕj�K4��S�X�⏦�T^�VG�-�Y��k��P�[j~}��j�s<�Hc)rc^�6H���B�D#��(���U���������`݇l�=m��vbc��!L����C�P�i�uݯܥ�[9ec�&M���k��f�X��!P���m��w�rأ!=��[�tm���8�%�C�����d�,�����EbN��}S�Zr��$tY|�6����n��:��k�	�`�ql��P$�.�T&r6�oQZ�%�"{��=ݙ����������!�ggZz�5��۰��ؒ��i���[�<�dUŠ��'���,jϛd����� `[)^"�c��Eq��I�P���Mpn�&�K~�liwb�>,�n�y72b�A�a�^���s��L}��K����`�n�n���vZ��!�eHk��;+�uǄE-m<yQ3��/��Rebu��oA�l�[��ݿ)�`�Q,/��xV��di6�5�m�&,|>}�]�k�>C��߅�wnc��-��נZ�R(r���8Ag�0�U�T����kQ�"V���U�*3�I���pI"W$F�9!S �R#i<�&�$��<D�SX�sYU�f(+X抌E(�%5(sͩQC�ԡ��Vd�y��@�O���(kTQAQ�D��u����TKK���:�X1��XU�
F�A�iiX�]M]TG;�J�T$21X��kEԪ�UkD5|�����d��S��p�E"�aC�HA��E���؊5�S�j�b��Ԩ�jD���j�*�:�`,?�
��<I�;(��QQ��(�DQF�b(�KlQEA�M0�?����yݗ���z�����
H���GK�����'�	/�3��,k�p�� ����72$��>��1�ǵ$��"�Љo� W�F��%E�[+�]���^�*��1�|���G���1������a��(i�}�L���)�7x�NmG���q.�1�@��L�D�R9��1�1�J�J�A���1t�a��bHu�*��Bn*[�9T�!,-0]'c�Zn��,0{���5]-��ͼ�s��ˈ�����<��S�KӞc��z��Nb�9���Ls�ck,Uv>e$�F\�D��X�4�¶(����t�q'�@�.<��:vX���k2Q�"���X�hIfz�S%��I��(�=9��N!�kN��4���B�a�M� ]�H�ӄ@C$H�iS�0�4d���e,&	5L����6���X�#)شѝq���J1�˩Dm8�<�/]�����F��Ĭq9�CS��}
�d,���p�5�H���%�O��-V��12����&������㥋�;�M&9��Q��d�z��E�L�B�ias=�&�x	ԣ7Ǡ�̥�C���炣�[2�C��k�9����b�b�G+M7�},b!���jE���՘a�%�ċ/!z�_ ����jщ�I1pZ< @ x�b$�%1(& U8�UE���o�=]BM�U��q���N0��Ҕuu�1C�A-�E+($O����P*sg�AO�_��<�2,���$��X� �9�����0-�+R��2~02 xq����d
�@<�����%��[��QU�k�,��X�[���T�d�~��R�T`����U�X��TSK%eI!�DAQ`�G�6���,�p:p�Ɣ9K�. �j�YԤD�TU���*J��R(%fH��dQLا�(���)Z�fA(TF}J��T�@R(N��0��d�*" ,XedU��C$R
E�
ʅ`,��2d<%QX�Y9�,�@9����QUN@�R$�E"2r@Xn��rr�~����HMO�	��RJ2k$�V!�-�U���,����/���Q���r,_��NJ[�;��[z�"�lQV}��H��V�$�		h

CV����FJ��f0����%6���"D� ��J��;�QE- (UE$�����(E��K����U@cl	P��-��A�A�!��2!�b�p�$�%`Q�T�J�!P�M�\������;��A��l�N��K�����}eg�ҡ� ��2�i����p��f���O����5�@j[�jOϮj�G��{�,�%&o�Ni��������T�N�yAÉ� @����	??�h�������P@:?_��[�=o�Q�}����}�:t��8�G���v��W�ϳ��-~W��%x��P����|r{�;>�� ���D�)|5��������C�e�語q� f ������?�IH~�1u�?���$��i3j��Q��}����N�#����B����,鿬�7�^���խ��`��'���Zk��d�_렧`�����v/���[��mz������g@��a'I#h|BNrK��x��h8�R�G� @  Q�.������v'�>��|\a�ې�����Y �S�g�3�f(7��,��,���q�X��|�d����o�-A����}�&u�NBS�;dd�UoGo��s5~T�Kn�3�]v��� ����.^(h|ع]vZ���o�|�x??Ƭ.���X��>T82��${._ �=�}�8g��kG`������}�j@����/��<��|��h���v�����<?��Y�j�m���qi���@����B ���+�!��!}VV4��{�=�x]���gkU��M,���{Ɩ���je�8�\�iT-����Z�c(�X 6�"�V����	i$�����UZ�mR@TH��b5F���U���*���dm��n010�����Ijе��0�c$D��-� ւ��!�Vն (Em�jX� �E��U�cce)*�ia%Q-�XV����ʀs�(����򌞴�g���4C���̜� ���Nn�9�fG�cc��[Cj�3�X
��� �(4�QI@�	�J��(� ��`d�B��3�RTD�Ag �@��3
��]a�,FE U �	XI��*�����>��0���*��&d�"��<�E��%���Af���@EI+�`�J���d�EQ#�*�P<ʨ�E���X|��$<��1D@P�@�
O0<��E�T��
���������,�aS�jd�E����`|Ç�X���E
21�	u
ȰYPQ&�0d�1LD�,Dc"��g�*,�3P�.PR!\�\RQL�G�E2��j�()-������9��!b�h������R�$���*�RC�,%1� �9��x(�)>�Q�1���*k]j��R�d�	��b� �H����_|1�k��Yci+3*�1AV

*(���*�$"�O�AO���a���T��%��+R�*5
��\JR�2�
���q9�]$0N�~����)Z�[lV�j)���B~!D>L��C�8�|�u�\�:�mC�rt��� T�mdS2X����mPR���aـ�3 �$� �Sy d�ME��´ii+k��S0Z �,�"��
I�@��3��ڒ�)��µN�P"��2�I˪�f���H��1EfB��3��d��� < O$���'��d��ʒ6Ѫ׋TUF*�h��V"�T+�	��@�-��3��'%[�촍��� "[UU-5��+X���*L��``O�O2@�$����>A`u�,��
��2DwԸ��4a`��Ĉ�GV�X���֕��$�>d�N<�.B�Y%jTVT*z�"���QQW�mVYP��Q��R�I�#�VBO$�|�B¤�0E��j���;�,�3��:�Q�UE�"�R�EQEX(�*�%�HbR�Ю��\!R	<�Y% `z�W�Bg����e\�Qb�h�3(��Z�"��1V[)�m��ś.���O~c;��TU:�=e����"�pŘ�Jҭ�M�4�*�4��I�,`R�Bĥ
���a$+�q3!�R��F ��R�����a*18�dE4���1PPST!�1CJ�U5UTM P4�%$�R���5H�4�AM)LQZhH��i��Mki�b�z�ڳ��R�pOOP{��lwI��h>�')�deʘ�=n �9��`�'%e�������q���N�l����^ǵ����������-�|��������x���[=��nw`��1�|������x�k�b�8�����s�����t�_�`��>=�z�߹hT�������tWGk=���e�2T(�s4�5z<Q��	n����r|^8�m���yR�|&g�ʇ��+�2b�P��ڪ�yHG5Lm���Ex8�f܎K�uq\4-��J8��}�~޽��^�����|�G�l~���~}�g����<4yW�L�߫�?'��=W ~�`Z���K�mxO������x�)I���M���?�އ��J���Y�nT�?�N+����Ħ��]�C(�cS��|s�}�V�ڴ ���z�"�;�*��^<�ݯDQ�1Gu��#MF�2���pX��m��Xax��g�ݚ{wYl�9.л�ˍ)+J��D�2�zg%���N�ZpH�[�j����ʋA�Xr(��©���A�[������I��e���]K�4�5�+Ὼ��&�[ �Nٯ�Ș�����<�X�d	PX���vMf���Qi��Pe��+|�6�n�n;(�ں�WU��P�p͚U�r�޺��1.��.�6�S�时k%,m�ʇ��d&�.�\;�	YV݀��-� ��3S�p%��6�2�f�lӐLo��ݸ	wt{�h�G��%/U&���q_EY�L%�̏R�zK�i	m��m�S9O/�r���`a���k9�M�xgi2V$�(CNF��DW�bT�6��\�5�vX^����>����{1�N�L:�.�æ�tF�Z���{ISHE�����yB��ݔK�.X�`��0@Eg4���Oa�.�sm�V]Yω�h��G9�ح���>�/N�h���C4��wl{O��M�=���F�b*��$}���ToB���X����E�}_`��Ծ=؆����B�dcՌ�#ˮ�/�{S�M2A�������,���(�%���2�ݖ��U��bo���EVl��;��M�eh�a&�%F@���$�g�oQƵ�NL��՟k�F�d	_��ϦJ�IZ.��3��=���b&����`[Env@6C�5���CG�&<���װFs�>}���U2�w��QWX7�J�3�����ˁ��h��R�e���q6�"bϵ6>�Y�Ո{��%�H|�l��	X>ė�,���~�|Y�N��a�=,V�S��� �@�� h@Ё�jЁ�K}��������7?�����-nO�Q0�k£������������`���X���������7c���q���a�E
'�#��k��<#C�v��z�>�?~�
��E�/W� Ƅ|Y�DcQ2�x����x+_��O�Si�䬩#�)?���X)D�;�����1��cR%�q�r<+�B˾�O����_%n)e�ٺ4*�L�\X¡��G�yh���B�8I��ȟw*8r������R��W+(\n%�K��f95$|��б�3!}ڄ(��Gk�Fa��F��PZ�nUV��A6PAc��9�c4e��#҃	��fX<�J�ԅKA2G]��(a4[�Ik����%«�H�����s�D�o6nc(z]K(�1C=.l��-ޥ*����!�3�BQH�U%P�p�� ��X��иTٖ`,�z����#r�ЧX
�S�1�2�U+A�3O@�
�=�T�1���e�4`8W��.,fͅ����G	pT��؜YH�5*(�;gD/L*(��d���P��z{� -կ%h ����8�T%�$z��o?���/�����S%�M�|��P����^��V+����ll6�)�'%�R�%j �*�R� �
J�ZF*(�*�d�,����P��� *1��RT��C���"��f���۞�6�F@!����f�����H�)�
 h��&Z��X�*1�\�hQ$]n	HR�I	*���<��{����o�8߳�~_�Q��ͳ����� 6� ��X����~�S���C�?�c~�?e�ۏ��(�?����	�g�xX��F��\�����~��q��{�^ߓ�Zx����u�r|����c�������/��Ol��������yا�����.%�3L~��V�
K�c�!E�@ �f�Ȉ�2dɆa���..�UQDDD #�L@�%)ƑlD�P�(��q�\a-�U�U���[*��)�)l+jFղ�Jڥ����}]�Y(u�Êuԍ-%�)�}���00,�	+z?W��Ϙ��w��g���sm�5z����AXb�;��(=9�����W��zΠU;��|�;�},��Qj�9!�7�k4P�4x1�G)��YV�T�UQ�j�o�f�#�����SE�8�x^uB��~_�(�3��tԶ!sG���   � H�zF�ܞ�X��z�'@��4(���VN��cE X
>�s�ă�z���2N�g��շB�������+s0gՆ��{V�M��<�k`��յ��]����YN��$%R��it轍\y�=��KǛNR�[{J�z|έ7�C߷��G�H�Ծ;�nZ�$g*��^��a�f��x�E�ƨ���%�\*Ά��N������0PB�4�i�e�Gv�R�k�*9� 3�dV�N���*��dcC%��)�m<$��c����ūF7��]��$_�	s,qd�L)a�u��i��
@����|��>t��G@�¦��J1��"<���q���,�\�K�wBҵh/[�;e1�S%�&GcE.�&�K�TV�%D�f���2W
�Z�� �B��ڂu^]�.��F4����:@�o7�e�ʐ\&����K��<\q�{�ϴ�<�
�D.�]ُ�,�H#1�G�\�L��;wiKŢb
b��F����RV�m�wBR��*�3���ضP]2����TD�X�?|�D�y���l��o-uI��h��z��k���iT����.H�|���st�~�X	:�w0�����P�T,�ї��1%pR��¸0̃nT�~�"�^��#j�]��ۆ���-���"%���"^�6��1���BGm�{M���$Q��u3���g�LvY�|h�Om�ƼES���4�(Q�a6��a�TjpGm�Ɋ��l�
&}g��F�h4`��V���"j���ؖYL�^�N�5+����T3�i�cJJu#A��
�A9y���T]�[z�x�w!�VArA�+��6Bn��j^�]�c�ە.:�KNѴI��4o�Wuky�i��yWv(��2�ץ�Et1� �V��   6�ՠ�ՠڴՠ�5~��_K���j�
+�dZH���O����ԗ�S���ӭ߷��qr}?�T�}�3����o�����Ϙǧe�ȉ&!K����b3[�x-,4�d�gu>��V���+�Q|!���W7�����gaW��)la�6�Ff�R ژUl��@Inx,�L�ly(�Pn����n�qfFс<�̹5�`˛R�P�ǪYu
�D�E��a(řjj��_8�8b�P�S�(/Va�93Á�� �
 �@���H�%�����,mF�u
Ӧ�x(�f(��X��"�^*`NfnH26�#^�V�Z��I�vq���M:��j���}VN1�l�� �Z��,��eP,%�&�F�pkŊ@��| Z�"}�'	�*������NT�P%�pTL\ۗ�As	�=X�º��<�j1>��%�c�Zd4��IT�x'JS��v�F�KU��[��M���H��(F�7b�߸�]�7H8���b1HY��'ʠ�=15C��j�`�h��Z/#����ߤ��Ã�l���F���q/Z�/D��/3Qʁ� m���R��Jb����&b�$�H�UH�!mTJ�2b�(RUFZX���4��Uc 2!É�D�R2�R�AT��JQBB�-(��-4PR!HR-�4�%Q4!IBR��IJ4�&�����
�(�&�&�%�L��*�ʃW���S��\�-��v��Z��a{�1�`P�ާ�|_�]�����'��_��t���=_�WY�.k�{>c6�x����q����i��[��O��~���@y�_�v(�Y�����=s�t�W_���QŔ���F�N*Ȇ�N KUE�D/}�ĵ(mK@�V�h �$��-һ���_�����W{��]7�v��	�v����׈;����;���������@��V�V��O0������Zйg�*����Gor)Ӧ����҅&2�wj�Â�z�TԹ&���_s����뷞�q�.m����
�	C
ȡx=�w^�݊���Y|�$�"A��̚q�t��w��H���OH��)K6���v-��)��:C]�����qUSwUK6�3O� { �z��D�����&挬NJ�E�%FuB��w]L*��9|�Lr��5�B�F�3ba��IK��]m8p�x_4S7�`p^ʤ���K~���4���ں�$B�-r��R$B�\�{m�YpF*C���΂��.��<�/,��?U:�W ��Uɇ�:�EB��4�H��꼢e��8�Y2^/T��)�-�]�%�r*�Y�qpj���̘�i.�0i-I��8�IxuɃ&��&�J`�	���ىﴥ�Z$��pT+��Y�L��h�Y%Ƿ��٨q�����q�PcU
)�0��~l�ذIM<[$���f���R]]ו�}�$��!2�QG�+)&p_�FP����['ۙ�@�6(̘�V�E^W,5ӣ$�� p;Vm�%uб���.�h��*P5�x�ō�ֿf 0+�R���B��.l�Baw29�Ji�v���2�$&k�#�f7,-�1!�1͕zL󊰈bJ%�^��2���9�+>����3R�w��;5���%}0B�DH�2M�޽�F]�Q�-{�jz��Z�ӑ��3)t�1��D����eU0�TEY�^i[F�E��+r��c	ä��}5S@z�d����s���9��OFVp�#js[҆�{�-yRa��;��CFKML�YZ]��o���n����*>ˆ��=�z��QR|f��#F$��A�+�=��fM����ދ6]IP�clR5�۲�K����H9r��a2�PC^$��{{D��/]���v<w\7#�q;�ZF����]W�Vq+���q�0)	^R��<-�\/���z��n���ɡِ�� 
���V�H��>�0q�P�����R��w��U��=��dg=�Is���Yn�h.��b��.�r�vB|�7K.,�s��cF�R�3�.�,�>������4�IM0AJ59�$Ru!g�Y���X��y�r���)$�D��u I�H��%W�%�gh�Te�R!5C-6ǀ�'Ɇ:9	��3b� qW���4Ӓ��txT-:J��MC���@�I'$�~�h5r5�˨���.�v룸���ŪF"�o8M�;���:��U%�BBaB�� �DEÆ�D�!a����~K�P^<A�H�R�ic�{�\�Pt%�g�,��!m ��n�b�m�	,�jq�[���Vɑ�ux8�^��$��0�xQ�1�w�9
E�"y��2e/*i��J�U*V�塣s����=߆�x��6������j��/�F���YqSU��x�����P��R�Ǭ�Y��Ã3l2f��l$*)������`pAT	1T%1��R�PTIK,TMe�TU08�*qb�s$P�	@��
b���B*Ph*���iL�`L@Q�8\*��=���Oj�]��~�$�����?���� �_�a�;��|���C�O�~n��{.��|G;���|�C?��:�����]�� �����p�yV�8���6�ÿ�_�Oߪ_����GS!�E��^����~[�k�o��[����:=�������O��\�Z�"!����w�gm�v<�)#�8����|��������5ҕP��e�bg�K�}�/�+��i������5o"�f������!�w�=|g�#�r:�YT���7|v�y�>@ s=���bZrG�W쏶/J@7��>��u췮jZ�Ȯ�#����f4�?_ev$
����\I��o�¾��El!�<����e0�3j�=$�Ԍ�	:&7�R���f1�YU����lӼ��=ᑂ��qIT�gHsvEK9N5��"٤%7ZɃY��-�j\��#4�'�������k/EDXr﫩�-���3p��i�4��0��E	��%3/l[���^�l�E���0T�6�m N1�ը�%z�؇�\����6{�-D��{�g#2�41_-��U5�˂�٧zk�oe�hb��-��C=�!�Ʈ��g(ʮ��z˯�ݘc������wI���J«tj�-
��l�����ќep	��YxZ�1��#:����d�5K�J�	[�j��f/j5��z�'k�}X��E��s$%cWi�v(��F��-(�f�~�I�W0vG�o>H�q�[}baݺ͓U�x2)4���Saѳb������GZ�y�Rq6(Ndl����5c��O\��k��$*��1��q�M��n���o!&���Ý�T=Zr6��57ly�����b�vǍ�&w�:ӗ#7!qc-޹��vN�O�^�a�I;1\N���v�$z�m�,�ڴ�,�,�'�`��rjLw9�K���3a��/71di\DU��~�Ӄ0��Q]kN����F�L �^|����ա=�7h�kq�0�=C.�U���#�0m�6��3i�F C%���hT��W�H[��ք�P�V��֋5���S��l�֦�׶,�xl�&�ح�pH�[+V�^���/��]y��ʺA�C�綝e���X[�d�(�,�����O6 YN��K�f�s�\�,pmk{w��jխ�Q�t}��?[��y�{����9:����(bC�󄤍۝m��|�l4������ Eߜ���_�O�x�<~�A@B�uVRQ�tr.���ivĉL,F�P�Y�p�WϮ�J4��E5f=\�0�13ԏ]�WHQ�u!I�͡4���(P�DB(F�Z�#!B��G�����&c��b��Hp
��k2��U��E�o����m�)*l�hV �����N8�IR,
�.5%�RP7�~_D����OX�:G'�8���/�C�qj{'�{z�.-�孀ĽH��k	
��5qB��AUjи�r�7Cu"�����*q�:�)$D-�R[�Z�n4
]&˦&����3s&� ��q|k��>���zV�RAd��Eh������t�����0�Q�x{�Y�������L\��'���S�==9v��S�/L��C[t��{|��S~(��j��C�ק��d$�@�/2z����BT3��[`�p\"3S�
���+��R$�6�i�X*	�`V"���EPDX �յ`T
D��$cZ	jX���7��P�A��lͤl�����P�
цV ����

�j���Ȍ{���^U���������xɔ�<�/���w�hrx�_��W�s^����q\1������X>G�3��0�������^��w����<���!�}oѽ{��_���y�rA�P��q�����(�Sw+�K����M�k�z��f�ލ�̌YW�f^�QڌTu\�*c%��cZ��6��yqu���>�z8����L�"���&&��I3�n;���]�2*�$v|���}Y:36��P�=�8���''��K]Kg��>�W3f��R,�����v�&�]]emrX3g����Fj�ɋ!�<�荹��1��TjX��A�����a�9}*�WQ�z��n\5�X���7.PVr�FNJ��L�F�+�A��-]],��-�^cq���汤�� �BL� @ ����;�9�r����t�^�iڇ����u����7i����Y��v
��`皋��[���f�@�����NWO�;��"�����|�Wμ�n�%��
�{�K�籹w��3\��<l�1�ŀ�j�W(����G�Γ3��Lr��a�Z�nf�˶�dd��.Wf��V�Is�U�z-�`{g}�uS0��pD�&�K�]gJ�n"�X;�jчY���w��^"sn�,�˫<�w��ې�v۝��.�t���W�+=a�a�-8�ǻ�AH6YS]A|lJWuɥS���%�9-�Sm�\�8��P,\�yv�������;�p�ńG�o�'�y.d�[�����uǊ��M�yd�8�#_�T:��]�����I��wdt���sl�5�*�o6��N�L���Sy+�v,x'���o�sR2Y0�c#�Ğ	���w+K�m|�� ��vl/&Z��#-h�{C�d�p}y�p��|V�l��rQ���`W�͝|���� &P^�%��6$_��ך�K����ٓRj�!$��� rZ1/Vio_0�Ԙ®�y3q�^\,j���Qj�ʂ��a	��$@��Ć�4>1���bP$L"ͱ܇�-:�")��4��%F2 ��,ߋ�Z�\˷y�G-W��C2�f���n�1�)�ˮ����|�@aZ�Ś�<�(�6ΞQ����&�V
�Fs��&,�
ykM�CT��]%,-�+`�$����y	2%5��zt�<*S�=1jv���f�<��0���=)��!��@_*�]�-�dQ\沁*A9�\P�V!>�؍	ujr���ED�"n�yf�j�^]�":'���9:ir�$U���lq�_e�h�Ӣ	��!ޅcf�M�+eY��1�%͚�q%�a�\سA�Ukv��2�D�30��e��&�;�e�s5Y�k��d������\kF�&`FBҠm���G��Ǧ�����n�����y��@dj�.��:ijQm����ՠLV� v�gmڈ"��b6�	�p�v$�0�]� �;���aw��I-3n�ky��5���H^oʠ�)ܼ+GXB�p,��ɖj���+�ڎ��,r��A�p�R{���,Tm��ѣ;L2l}���"i� �V&�����|p����}��0kP���A�����A㥝�ڝ	��<�9�E=�L��0t��r�H��G��5�]�^?��{��k��? ��.x�C��_�'�o�m�/\|o���*�5�s�#��ȩ�م�)a!呑F�&]t�R6f��`�ى"�-Ap%�,�j�3a"%i�[5�x��hv��"v!&A��	�e@M��E�	�0x	8�Hc&Wie�j<��
,��(�%�(�?��e�,r<�}2w��R�X�9�L�D?��-�T��EeJ	$��(���d���\�Qm�"��TF`=ޤ�6�l�V��id�
�L�#*!�K�V(�'0��t�$�-�R�2V"�i�h"��iml-����lnXO����W��~C��\����]�O^����}!��+�~������<���|?��^=~�zg���[��=��!�>�g�<�k��'��Og��?�츿U�t��Z�h=�y�9���'�?׿������d�e����gp�+��\�{��цL�+�����AE*��S1ʔ��i�]�E�d��볁� ��x��.����\�$ڜX&d��6"�T����Ͷ%A��ǩFuXY�yU�gv�4M�/i���8}�2�j��f�ZG3H�֖�2o��Yf��\��s��|���=,Ƈ1yV|����)ۃuX�E�J�+�Uչ5�T-]���vr��2��ۛ���;�W��I������Xm-R3��W�MU���y�E�*|V+fm�Gح��y����Y�^U̹��"ʝ͸�=s�
���ѢO�L��5��U�dw#Ã�T�̭}�f��	�����̈́1�TU�ɨ[��.�[^wn�]Z{	�=�S���ؖ���F��O���i���������-���������/��<��YS;~C��{P�M�x�ی��� J=WTd�L���[��{���Ө���Vb�Qߞc��^����wGw�q��"��G@ S��([�L-����C.fa۶Źb���s���"I��"z���5Y�t��E7t\ЮgU3Zn�rx��ew�y���;�κM���6��F��N�$eĤ�t�5��"w!�ޖ#5i�&���dXA~[��8����ٛ�i����q���l୤H{�6.�i&�3�B���=�.8�N�^�n�<�e�b�(=��M�ˉm'>���p��a�)�V!����}&�Z)/TFm�}-���/�n^�AO�Iz3[�7L�I$&4�\�v�uc�M���YUM���s�!4Q]�m��M��[���l��mM�S�X���ͅ�z�Љ\���!K�p,�Wߢ�5ސ���5���J(��q�3��焜�k.�1j�Z���K����B7��M�Хu]n�}f��GD�MP��S+w�R�B�E��,5H�Q��@�[J�wt�Jk��&�V��2M�P��$�ͷ��X&R1�s��K�1�9c�����fdm(��g��N���A��hY�������Wv�g�L�MrZӡ=��1r��Dw�PԢf('>��^�j�7ֱ�NX��/R�!*+����~d�L,���k]�ʿ�	q�E-`5����. ���h,�Z�����TY�Lds�	ێ�)e��V�ނ�g@v
�-3�mꮎ�щ�!vE�$ŎXF�{nR�xw�}B�NrGь���-�a��[�ձɹ<����7�լ��U4pώ G'����|�$�L����]V��tK�Ӫ͌,�8f{�*T��1H�洡3kJ�&o>D�E|��`�,�t��9Y�Ä���!"��,%�%�G�Mӑ�Kz�6<P��g�8-v'6�*J��1x2�]�h���p�a7va��A{1F�I{`M���4���D3�c N��D#��I&�$ ��b]דv�#w	�sc�ʩ�Q�K�yAy^��D2E
�'��g��,t�ː���+��w�=�,V���"���8�o���.��{�ai�e���B=o�H4���t���??^*�钩�X����V$�BG�E�ޒE	@w@YK%0?	�@�(h�c��3�E�N���i�$]$Ъ�����@��ewBjm*�"��*۫H(�6;�;`t�T��Yj8"�� TF0Cyp�|��qc�sݺ4f�<&2��/O���%b>^N^<��}1�3,���D���ꌋ��GEU,KmX�	(��Ȃ�A���cl���zQ�D�[ �d����*V@Y"�IU����N� @� �'�n~����?c��I�3�t��G��9~��p>��y^-�|���s~Cԗ�w�?��:�G�v^?��#�f�>���������Ӓ�G���d���n+Z��x�"1���f�����"`�f
(( ��`&!�"�"&"��" ����"I���J���60�Q�� ڌ�����S  ����9�~���^dMt�s���F_FQ�Hn�{�����7��@	E��@ ��   ��;�+�T����������  ;"�S"p�j,q�u>'�vkŹs���k����v&��x�;��v�e�c��sEh���h��m�:�N��,��O���W&n�aH�!>'D�B@��z2[9Z>��Y��6ŬA�s"Qp�{�v�K�|��X��]�
H`K.�	m\�=J�G�)� �ˠe��ə�������@��L
&�Oh�a�h2�e��P�U0Z*@����-�-߮<����6ֲҒ6O��͊>;h��XW!�5���}�g��igc�βe��U̅����шdn+a�*�R���'�:�4�k$y�c:W�sV�7.ކ�y��>�Y#%����W�+zp�r*-sVf!7-'$�a�C5�����U{'0Gce�fI='�R�ܸ<ZT�o�-]Y�/,J�J�%�z�b�$,0El:(I#�A�HRN����']8���T'�{5�(^LP��՚�dR`�KɈ�d>���$$)2�{�I�ډ	�T��

@�!xT��z�5�KړTr�'���<j(��HۗM~�C��2�2]�8��v��zU�K-�Cn(5�1�#��	(k���F]6�_9IΪ7�j�C�;M7���Ma<���cO�IqL�Q^��Ҟp_������&�� f��l�i�&�E+�7y��������~!�o1�C	pF��V-U�����H���ZЉZ��ʸn��B���=
���o�~}G���_
��I��L1�oj9�뚣#��))���ɉH�J�ؕ�Q�{��Ҭ�և1 ���L5}b�˞�c�VgV���o�*��Y�ы�+�n��B�(L�f�N�܋S&�N|�\i�X�-����Ԍh��j�N�/�~��L̷X��&1����S�m wY1]碫`���U7�NF,0��'-�Z���P��Z�<g��<�o�tz:N�s���r���?��r���u���
�v	J!eXz��X�E<�X#�(�Fg�9d��]���ZN�W��)�Xo���l�B�5�#�w׎���8x礓�:�o~W���o���D�^y߼;���M��|v��m���˪A^3��o�9���}�m#����X�p�NݩX��im�ϲ=�w��u���Q�,������âwG�ϧv���Ǐ�9��ÿ��
i6;Ӕ��0��V��t��n�/}�nq�K�`�C��Ã��0 �H
���$�����s"l�e
A�N⃴rjkx&&	�lZF�J)mkH�`�p��J�*�)�-�bk���	��.0t�↴ |��{?7��9�GO��h�|i��K��O�g����{���Jy_/�G���{��{�S�}g������o�������������_��/�<W�����tt\��w� ��_�~����g�����Q�f���D�mkH��\*�k+��t\UOj�����5�$��p}�3��jc�����Ʀr��L�wV��.K�]��l`�#s�[쾝�MR�;��)Ӆ�d�oa���M\`���yx{v�d�(�	�rgt��֠r�}��TNz�F�vI���o=�����.�b>�T�1R+rOA�gf�ܔ��ٺ��5�Ĵ1HF6�r-�(��c	�9�I�λ#Oi�g2�Dc���sӗ�ݣ�߹�V�������Pr�����A�_PBcb����3 �V�������-oZ���7��d�)���WY�ѵz�j93yN�F����:�Eȕ�u��R����͛�%�V8d��/ܡB��b�i6"��Ω͚�r%�FhA���B�DD]/,#BE�B�,���E��Nx�����M�d��2�n�rfuadU'�$Y��y��2�p�5Xqۓ��F�Q�f�^.����wX�5{�a�A����Ό����CR�N3�X�i�����]�&�]gd�e�LOPG_<b�j�����Uy��-3��n{QR2������W[��jQI4`hUi�����Vk.j���WWr��ҷ
mi��5qSg6�x���ک�1���D���DC��ڬUs�@�{5]"i�z�p֬�9J���I�
�Dl/������^���x�T��kt���RJ�DH�ːZܹw^P�����c+zM.�'�*f�k]�j�����d�DkP#UNF=se�=�_��p��ױYs�إH�˞������)�A���iLS�n�'Qp��3��q[q���n�-Jښ͜��=��fV�(�P���NM�I�@Q� ����Vm�K�M�Kj"�殪�W~����>�U���z�9=���B�w;
~��+�&	ݮ�;����h��U�>J�6..8ӎ$u�a���x,�����s6�NV�	���[�4^b�Rst�qȘ�������0��i�5�ن�X��$�n����7���ݱY2ާ��q<[�]�|�ڃ�Q�8q�DD�uKkj�EmL����.�2��=�y�w���������Yy7B�m=u��ۭ�y!�V�ӅJ�v�NF�U;�'�S��+��Yo�D�{������5���a�l�J7 t��������9=W��׷�ʷm�#\$t�tR7S�+o�a�V�a���C{*��n+"*Q��X�nz��nv9�^4���[��I<3�8佝u��:+�F�j��Tma"2F���8&j:%�US*#j�0�H�]<7j���õ�{+nc����A�νH�w'���y[��ݻ��=�c�����z����F�S�7�gTP�(��/C��W;BgҌ�0b�\`�󳫫yd����DW,�~��n����
��q���//��f9gD�zc�����W���*��:t^�ۄ��"	�n�N��]�����"������OGe��,��yd�kr-ģ�S&�0a�!��f��P*j8]��u��]K�/8�4��TE�����)Y�38rx,�0so�'e��7�ʏs&�b{2K��"&���d^Dļ�:�ѣ^s��4������0�l)���X�ES��I�P��u���̼�&��6�7�Nk��kg:�=4=�Qr��~���세FN;
����6�-����;Y�*s(c�Xqf�MV��쫩�֤G�f����8�:���W]*{MI���FUI�fUt���ܭ�&4��H��`��nٳr�n�S\n 0C5��ɑ�iO(�H,[�4�{sZ�{;��9����H����Û�����IX�7]���n�2��� ��v�V�3g&g�n�!.�{g2� �2�,��@�#O;�]�>�kQ�9���Rz�B��W���J����ѝ�ۛ���z���xlS��:l�K(�a�t�V����J�
�M��vCȫWTh-ڭ����Iqx���k��fd���[�w�kQNՋy�f$���iϙ6MkWB�F��ڢ�;�Ck���3�q��4�ݸ�de�8D�����ۖ4�M�hÌக�E���3~�Ej�r�PT�Q��6}�채��t��rڴ�3�"Nݧ�]�z�.|�g�w����K��j��.���l5���§e����R�Z���j洄c���g)Pw
*l���� tj�g��nf�!)�Q]�����gVg0FǓ�����p���Fw0��P��Q��9iDS��ԣ��vԪ+��-�
)t���軧��[PJc2��uYp�&5Ƃ{l��[0:[vr�y��]lEi5�,��ݙ�S.6q��|�zWf.�ᶋ�)[�*������Ѵ��4"Tn���unޜ"����I��P����+.5;�:���Qޞ�3.�$vL�b�TulG���=ۋ�e�F�b=s��'6eιf���x�
53�.�l����%I]���|�N��V��9Y��#���wQy�@���۲��]S��t���<G@踢���95XLu��$�G:ѝ����f��)��#�:�X3���%&2K�Ϸ�c�I�v���
����f�����c`ga�W�>JsL�݃8U�d멠o;^(�1lɵ�nġϯ��u~Z��{3��8P�ld��}=��������yq
����Ҭ�uE\�]�"Zu�}�-�u�y>�Էf\F�����+#hr��h�9�8������^\�i�=����9��S⁷۳C'E����܌���kb�4BC54����̧�=��P,ڙy��w��Wi�J�nt
�\�d���1]�c�2�k:�ŪZx�S
�{s�'Dl�	u�F��n���Q�b�yKP0�4A�B]�V�VKy�lڙ>fn�4�:�U�;;Q9�Z�UZ�PC��MG9��N��WB�˾���3uՃ�#��x5�Nб=Ӫy�Ke��̢ιT ڐ��1S�E2�y[���E���UR��@�d]/��ц��3"o6*q��u�v��Y:�`�	�@۔6n�Vo_e�ڊ�gg�[������*GMF��2��9[0���o�t+�b��kf##aj��4�V��#�nkD�;��9��3c����鋍�".uf�̗�V�Ҡ��*Xyp����^Un��f�E�n��ޅg 3Up݇=
za���uj��܉¯��q���T������ƶ8����̈́$e�nzs��`�U��/15z�6 cyj�٭�b�.'4a+�EN���.���{H�5�q7>�c��՞�ϱ�U���r��W�2��Qk���=���Λ�hfu�8��)py�4:�1�1�*�ëK��Ь�Ή�N"�]�גhWS���t�A�9:�r��@`.7.��jv�l�KQ��P�x��W^�5��>�3�l�K۩܎\Ch����L�p�y��sݲ�4�i�!�s3ؒ�������!N����j��Q��(m'����`�W�63]D�	M�v�ѐ�{��u!�A��5�����֮�F��E.ׇ�d�;�W-�d�W�]�Lcu�rI��(����j# ��B9Rs��}��x��.���9]:��+E�5��e���j�ˮ�W����3	�H��G>03T�F��sgGc"ZW���A'��/VW�������9���f]pu��(��UFb\�
٧Y�¢o����S�$.�jF6������t;7Wb����s�ȓz��J�����&_U$擘���I��4g��Z�{Ѷ�e����3�g=��R"���5z��v��2�����[zFɸ���ZnA���r�d��q��XQ�8a���ʓm=Z2�;�xvu�bFL������]�WZ�gj���f����/��N�B,�ͻ����򧦶�t7�
��"1x�OD���k^-/�u�:�w�fm�[:����l3�\��5t�ya%Lƻ�g��^F*��婣�����H�O�N�9�;�Ș��n
癐-�$��+ؽ}�����ȉʍ��&)Z�}wP8DV7����;N�ˉ>�깘�̘�P�ғ�O��:�v�ᚩ!l���{�H����Ь��z��
2��a͍>�h�>׺rw4Vמ�7��Ɂ����^���I�вw3�������SX�Vtn�w�v�d���\y�ba/v�����Χ�]�7���&�D�2r:V�욝��v�w;�wT.���k9�]|����PFۍ��u�xxt��:�NUR%͋�
��H�E�':�ъq���&�g�b�K�ŕ5̤��]c�����:3'S��fd):ڌ�W��"�33[ǳ�<�g*��Z)�]QPU�c(�=��]�v�(�X6���)�l����lveCz�2���W��i��|��ԓ	v�|���E�xq�2lF	�9����L>���\�
]V:6"u��{5
�W�IO+ gK�b.����mf�Eī��޲���L�!�$�b�	權�hL�_3�;�疽�W�f��N�[Nz���J��87w`�<�# �Y*n��#��dޛ�YD�r�+�UݣN���;.��o�f_����r�8��c+�:��#p��}3�j632�s�1��8I�ޡZ��Ki�ٮz��R,��t_��q ���u�t�n���kk�t8Vlm�C��e�B���)�ƈ�}4�a8SF�<�8���w�A������ud�dh&7#�R����wfeY{�䒔��1S0����b6s����{�2$[;�����V�O- ��Vbn���22��*b�ʕe�����.��LUN]1u��`�:��29swsuZ/{P$� ��x��{�3�7e���8^�Q�5��E*ڻ�ʨ�a+�����L�Z1,+9/��:�U����
�ge�Y��
5t�{rrv�%�M�,o{F�҄xYyi�2�L�n�������x��m%�٠`L*[���_M���n;̉��q��;:F���@͢l��E޸K���B��($�y�+n
��8�]�����6�M�ֳ!�FN�O4��e��#����/6b���	�qWюsue��-h�B��Q+��L�N�u�)�ކ�E<��l`�3n��ժg�BƠ�����I������;����iQ9.EH=�2����"�H89m%uO:;8���gWW���vO	�b��{}�{m\md�7R�xlYw5�4�FNh�P{ڏlK��z�����m@λ;q������V�n\DMNoK�T���ʩ��B��A�}�H�wZ7��+1�=W¨��kQ�7F����]9C2r�dkۺ�����}[D͞]:�,�7y�2��*��.U���(p���)�4�-�eթ�{uC:�{4Jǆh͡uԝB����y�<��������Ȋ�L҆�"��C�wve��.�v'��L�kS�Q}Z�ٙ/�i�GH6'$U�Nf�V��OM�1��̂�,�Op1'��sw�Y��#b�8����1���`d�����bJi��%ke����Vm5QII
�#T�P$J�b�&��Ah����#�!)@U+�LDB��V`�d�Q��Bq�l´Jʐ�
�R�PX)�jI+
�b��B�@�JD��ZP��Ć
�EF-F*����XEQDDb�E��+mlj�P,J""��Q`���%dDH��QB�B
B�d�+
�V)X
dkaYY+
ŁQH�(�E�*��H)P��E	D��"$�*�R!P�
 �ImQ�� m��T�R�)D���@��J% P�0,*-E�k��%H�V�J�h1���`iJ����D��b��DkH�d�� ,�PXVJ�VX��B(,+
�Vb���(()
��k%H�RV[i �+h)�h����"��X�IP��Fڀ�*k �-�,��R�Ԝ`ڑ�#eM�l-���I�+�$��G 'E��}���,ݛ����<���Ǿ�_�:=���ˤ� ;v�W����C�L�!�9��y���LcP�~,�v����-)	��ѐ�}��v�s��+���W�G3�d��Z"�[ k��j�/
�}�d�&.�r�G�����K��N�F�7(:��ʑEitǡ�Z	M���a��d����bq���P�uY��N
,>>�:5�X\����[�1m��/�h�]-����,#�1z|op��t-61*��!��(L($M�3j�φT_�f
Δ�+��/�.WKƹp]x�����t���9<ɷm�Nq/�^�9X�2�\6��{5(o�����w�aKZcz(���۰}7�Q�ԣ�$���y���#7b�z�x�`S�SfGd0
�-�]8�j��l��KHr�4m�Ŏ�ҿaG�G�D�E�6����خ`WI�dBcF���^���v�^Y�������R�P%�����Z�S�7�E�6Ly
��AD��h ��	�ce��!	���`ʭۈ^[��@�ɹNdL�`i����,��q����M}�5䡍:E<��ڞ,wvL��.���4	�ye������Y��h1��tVt�&g��%�俤�爔�7�`��&C���6���ڳ%$�Kfӥ۫��$�a��{5{l�Ӣ�]&�۷��'z����8�m��@S%rP\ˊOV}f�͸�I/���q�{�klYv4�t4�+$b���Q]�Z�ݣ޿m�˚�0�+cz��J��"���[ۉ����%e�]yd��Do�|l���[\/������ԉ�ݷ���gB��0�eߞL۳�So��A/d��E��cF�(�+�t��>���Ғ����ν��أ��iѤ:+��˭ �`���ս�][�j�N;���$Q'��h��+��򕶨6�d��Jd�6[���W��Y@Qp�u�$�Kd;�&�e�^S��D�!1��71	)9��XRw����i�{<"ML�Vs!Z��.�"�%��h���X��P��0%�s�0q
/�`��|����	��(
2E�Ƞ���Ǡ0˨�n��I3TAy%HYb�U���i��i2�ֵ���_��t���W�B-q��v�����p��{5ӈ3ۊ�����-4�?9P�A����)[G�ϟYQ�oD�g
,x��yr�l����.�.X�(|���8�|����3�k��3�;��#�p��Տ��I[^p�ˏ=s��Z5s<FFb�*�x�� ?٘��C���I)���QXHK\�N�+b��$KIU� �Hf��DE%-bq&aW����ܷ���|���y������%{����>�������4�'�r�q?S��x|/u黏u�{�K������zM�_����s~�{}��������*�a�rA{�a\��X �:��9�����������y������>����y��C"@Hc�#;�"�Nt���P �D�F�=�����/I�I���\�t��U�zb�<�4���L ��E�D�O �����U  �  �p%N;��j��$�0��GX*�j�H2�$��1�b�ԗ�̥v%tiuz��Z՝b�	?Z���3�j�n��6L�^n���{�h�e#V��QXW��z�(���;\��ܙ6�-�J�U��t>��Cy���ζ3o'L�Q#Vw\�6�
c	��+ �]6�w0�x���c.���x�4�b�Q�8��0Z(�sE��z�x�c�&"��2�ӝd�P�⹝A/����\��}���n��V�±��"7��\����fv�$����G(g�@��C��|�$+d�d���T���[�^�4��[Fu�k�0yj?y��.줄��8�h �L�1^�&��vk3ٸ-�c-�ر�V��*Q���p��d���ʩ��(B��cJ���#"���P왘�[� �L)������I�����Ѥ��:�w�~�hdwc+��&a���V< �M��$���ᤉ�ё���j��֋z6"�/��,�ݖ|ƜH�2f���M��̩oA���m:�M�X3n]������%6��C��sJ��br�u9��O�6���ˈ�"Q�Y=��;�ѵmȔ!�)�!�;$KTi5C{��n�i��-��~-B��^�����7*���fc�,�6,����Ϯ�ӃX�2x�,�.2�ƅ.̐��4�p�O��VL����3^�	�N �i[�V�r��S�	kbn"�ÛFXt\xE��o�1�ޔ��80ѶY��z5lN�z�k���"`Ip ��W_(��^��.Coo,@�5S��F�ӶQ��4�Ipgq�ӫ�H��-i�{K�36��pl�'�t��������6L�ls$��Ȏ���h�̎�wo_�e�����6<wP�}���Ԁ  � �p� :�����)a�0��|A�Ԛ?Vw�C�G�$�M�܏LBd�ȊJ8��ESľ��ZN�d��Vl���}�1&^2�&Ş0��5	�s�-��V�<�y�M8p=5a��C��X$��i&<�.�c�r�D�γ�x�ʻx��i���5��R�����h��g9R�=�q�%a[��kSK�5����d�����teٯ���0� � �p�����N�����iV%���eZ����`�MT��2ME����-V����&��d���lͱ��j+>����&�����aĢ�� �I(�1VEl�P�����{�hȢ���c�v���|oY���\�e����y���G̽�%�߂V��;t�s��g�l�޹Oe�v������O��k�s�����|�Z  ��Z�K��G%<w����9�a(��(��p����=�����e�l�2�v��saմ�i��v�iil��hJ�Η�6�%C�mGS�T�$-���$:+%�1H�S��C�(*�ev�!�?��vk�ց3�f)�ΐz����R׀<���]����T��G�k\!�1M -���]����� c��� v��S�0	(���ګ_\�+�SH�3V���H��a�$�M&;��}�S��\fە�����G ��zϢ��o���?S��^�(���y��~��Zߛ�������7)�{������K��_��K�� �^��9j�)s�s�hUqAar���}$���S+�b�`�ej�dhdi5j��?9�ޅ6_�?ƶ�?<;��������pfj�I0�F�N���kM�J��^ZRiV��&���(�����YC��1d�U�H�6�B��h��phrd���w$H\J֫�
����H�Y�`��)�󉝠�<���(f$iI$I�$���QIM4W%b�#&`fH� �PlM�bڤmM��l��i�)ZE
i�h�
B�C���<�v������tߛ|��c�q[�~��|���s���j�o�����y/q���^[����q�<���
z!u����YF|#�2�m��D�M.Û����?�_�)�Kg������ g���>olYʅH�9��uf�W����K1v-�t͵��h������y�_�������O��?�� ��?��W�蘆dg�əV�.*N3��0h6� @V��q�{^Ց:��������r���]Y����x�ۄ�]7O��u����4�'��8?�<���z���}[����_����W�������Q]���!A$�F@�f�搐���fc�����|}~=�S�Ͻ����eQ+���Я��|��=�������	�D���4rQL���[ũ�|�x��Xl��1�p��Ad�U"�ev�R�q����%g��%��JⰧ���e|Oտ�������s����V�%�G��6��(-I'�"��/�B��%h������1|��~^���py�2�C�rhP�2 @��G����=�3!G�d8d �#��_^����},u͞�J����#EF��ҳ����J���G��yC���{�a��s�|?O6�K��g�o��F�'\�m�Z����dV�V*fԜ�M�=����UQ���~v>�Է�B�ow�Tɰ� ��ϩv��"���5�����I���E�=�/�D\M�ڴ�Au�4}*֮���Q���/�~����5�mCۧ!��쬢P���rVV���^'*C�{:J(��t$��k�Ud�I&q��ʁ��� i�B�ej⼙��Đf��Y�0�d��_�_�8��i�w��b���ǯ%M5�֊�Z�0�Aڝ���X�\��n��P�G������4V�vB�BU���0m���w��$"=lf���s/3���&%C��ds��D`"U3���;�@��#�Y�s��:Щ�Jh�h� ��6�S����e���b#� ��˯��&���4I�/�� �u]�2�izT���2l^�'�J��������a�^�/���9�n�Had��͎�ϛr+#�����)B-������B� �:ٌsX�ҁ��(��u������oI�X��r����`�zr��悓,�>F���p&k�Z�u��4��G�=o�PN֙����7�Y9�bE����W���w�K���Z�>H�O��Rr��ڠ�R�E���OIP�4�,*��\dd��#�%p��*F��ZJG���L�{��!52�iJ���
'g3�tCH��X��8��D"��8���Nn+c3��erY����o��~�������FB'giQ�˳}a��
8�8�N�-r�����;6Mi4�f�9� �E'ڗ+Vur[-2˙��@��35t�`$v18�h&��dqG'sy0�rCx?Q�58
�4C=�G�����23�JI����&I�����\���X1���0`�$e9͓]�Fb�cMNh��F�r����6\,q����mU�'g S�"�4D{����r�HU���	� H6bv$��t:�Ϊ�j,�܇�� ��:�,��)�l�g�Y��i���TmQ�B`�#!�2倃3�l�K
,�������|*����ƌ��^3J"��
4Y
֔|��2g�͖%����� ����?���I��aѱ3vB�b2X��a�K��6�I3]d.tt'�LEXBF�D�.�$^��>C�Lq4�4L6p���#!���Sѫr+��>���!��<���k)�D��������"�H$���"g֊q�34r�p�3�ɦ�v���pA2�Q,�YBb�#���ΎZ�� ,3�22�;52/����?tt��^�2O���eYTMW(�p� 2;Y�f�Ey׌E+uS�[͂�Q�(&�AZ��a����Q.)QX�+�D����	�I��DF���X�oc��� ��x�.n���Ϸ���h�������¼��]�vy
^ ����	VPX%�q8^[g�q���C��ci�}2L!� ���O��i�|�`'UD����e'�����O�A9=��!GG��O��"�#HI����<��0CVWdy���	�1T��kݮ�fQ�����$����cUS�R�����s��J �OKg%*dL�ɝ����,̑�ŭyD�2g#�E%v�d#��f �)����v�9���9�6��u<p��lC)~�@�p%�|���Ҽ�e8���#���Y��WFcD"�{�!�Q�I��@�������W�N�#�u�1����lL"4=���L��]�p6C��bR4 f��*C��u��7�t��B�E��
�����Bԁ���B(�����5�N&h�"�13�x�E@3%�{U�����9��؀��c�P	L䑓�3#2�߼��7,i�Lp0{%�9�g��B"��f�O��f�D0|�l ��!-:��zl�RA_�D|G��>�P�4���"�F@�b�5�@�dj(D�l��h�6t��hFez��SaCD&�f5��@�����R20:h�J�s��e0��D��@��L���#a/�x�?����R/�<6ZP�Ȃ�
G�0�g����h46�H�1�P+�]�F��`	�L�a8Q�)p�s����Ch�]+��d�E#c�:��M��t��d�AkD���C0*����9"" �NaWS��$�ټI�����������H����i$R�àmh�f��$�w4���0Fo�c����`�C�?>o�<1'�~������>��#$ �hi�%j�U5M�a$���b���
_b��(P#/���6h�R���L��fG�֑ń�?d{I4m�����9��(O�6ݫP��@�h�ba*fT/P�	 Կ�~�Q@�nܗ^(g����;P}�]:�O��s?����U�g �}�E}��П�Hk�4����M�;>~�}j��`�X��_��c6��3�*Ҋ9�%ϴ�"�7DSS��A;MMa��q8	�2�T�$C� �(;a�{ĵ��p�&�,5nnP�� �	j���h��_�h��v���3+�e"�����F��t��-ܞ�����w�b?N�)�ُ�2!�� �/\��]**�eB�#������_�\6ˈ���"�f%�4���! �4�P�R)���	�����?X�V���!��r����kn�YW�q�{����L�#�������#&���?�o�����z�k2���~���B4A��F8��SR)�[b����r�#�7E���E ���&ߧD/⵴��}M�]�Q��浮��Z�S"��Ia�)FP�	/)G�&�'��t���M( ��4�'�Dõʑ���D6���������JP�l�	�{�&�3�T~~ע}�2���_yb�)����l�]8ODmh��{'�Mt�F�י(ʡ#�s�BɰYœ;j�R�`������fDE�� ������9U�<+Q��?t>�ǭw�.�`ב��Sr��E��������tKIn���ػT&ՔX6k����o������!~S�P�)Kk?עN��o?7++y�4=joR�JPAP�6M:$GS�)Y���{��ӣG`��� c[�'�Rj37�����I&��4��b�
5��Bj�'6��x�f/J�Tb�JR��VgGzgr�028�����A2�+�Ոb��`?@��C�0UrY@ @�/7�<-�{:H�̜�g�:YV�C-Z�f�f��l�
�f�b��l�,%_���9~���#I��F�t_�(ή���n�D��d؏���M}��X����xdB����Moy��P4��������z>lz]�`�9i�����,�̕*v{/-��8gz��dN/��`v9[9g�M*$h��Jp�g^9�1�Id&�:�3C��~/6�����O)EP�T��[�H�@������qcA~��sέ	���,N!fU�M�M.T���`�$�1[D,��"�ew�W�0�������Ns���L��X�w���XD���(��#)դn�x��p(��R`�pXу�Q��K$:�#)��7�O��Ȅ�'߇��]YVE�Md�ғ��"�V�)�V%(�
�\�)�R4	��@-�
գ��]�	H�L��D:�J����ۢ���#G���H���g��$���g	�i��{ V#{�;���g;2�0�� �o�X������w=1��Si�h^x�Ⳬ&�Hx5���v����+ZS��Ƞ�q'���Ԍ�����W�.��*�$Wy@�o�'�lbK% iiC���Ǥ�Q	���ưA�Q���Af��b��ࢡ$�p�U�#"�=�бw��Ny%沁X�h�G�O'�Ҍ0�c	l�q�q�S���S"�d/1)W&���°��u��m�>�!�}��w�ٺ@���.��l�ER$39"`T�xJ��W���?>�!�e@����13L��*%�"WG81�:��21b����� !7��L��� ��%g��!�U�����!g��y�i��ILB��)P�Vy"�ڶ}<��׃<�_�Z=�G�}eq����:*�<y^�iv�T�ѣUcJG��Mc7�g��Y���T�5dº�{�t��r%A��A�#cZ�`q���mqa����.V� �#��F92Nz*v�ggP�� ��s�G����͜�� ["kUZ����}�[��LP�U5b���α�"�$�<^-�"3 �]���(�6�rA��,�ik��!gAV�,��DNե��'�%�N}I�`�9������a�N�Z9�@I�x6jbfw�R1���RKр�h3_Q���ߑ��� ��Z8WϾl��=Z'LI����!���'�JGM2������k�����4�ivYQ�'9��T��gZ�jHD9��"Z"sh�:��S�Q�9�d(��_tgY�ʆ(��ʷ_���Y���4W���=�Y�6�]�e~����O����BB�a���9VH+t��x8����it@tC��xBKH��NP3�Q��b�s����)�s`��S�͡ "�m��˜yȜD����F��\�a0���Vl�V2�C��� �a
t��H��긆��D$�iI�E�%,���vʴ�3�����˟/�y�c��QT�s���6������Q(@��)S�0t)��|Q#s�����C�����.w���rw�S,���s�+H9������}�#���ˣ�����`��+��D�hi|�Y	1Mr͊�8d�S�LwI2B�bY��c���R���N���2���04�H0z��$�7��z��Ŧ) ��k<JG�K=���F��I�<aD��ZA��ʩ"��%xCIbA�^(&�	�&Љ�gc|����t�#���},���W���A��R3�2�#Bt���`������C9��IE��)�Q�
x����gm:�gJU���j�=��:�0�����������%l�I�4���	0C�l8�|&`��}��e�! �!��c*8@yB�29���qQs���B�::_�������%45l̮`�3Y�(HRr!g���U�*�L��s�Jǉ!�N��T1C�8���ԉ�I��SC{�LH�J�@�X
�dO��e�ǿ6y���v�\1�>�|�^}X���/��5�]����4��|E������O�ez������0ՌX�0�bh��D����Fu�E#
p���s�C(�4CD�S�?7���`�Q5=qU2�	#���l`�GT@
�:C�X� d�B���N��&��l����*`���B3TD �S�� `���z80���!�ݘ$!�~8jN�I����y���r��H?�we��	��e�6E��%.yx߿F�rXf~����?}���B���?X<�df"����P�v��Kɲ|��݃jP��k��
>(�Rύ�s�����&� �B�:�j�#5ɂ}X�%#	{�G�`$B����ǆRJݑ��%!!�J |�߾����:K%!߾pD�w�b�� �������$A!y�LzI�Ǆ�2�9����p5Q��29��A����ߴ7O�"R(	�I �VDğ�͘?�����6:�~�����3��4Ke����h��W�$~ĉ3h�?9>�_�VR$-�<�@H��J ?9�Ǫ]Ų1(�}�uVN��	Y�K�R�%���$Ǘ߂�~��
u?bE��
	-�z`��+v\/��B���f	�vMM+Bfl�X�LׄIG�cUi���;����-$SbDu2>�zF�4���ٝ��x$��)�0���_��5��y�T�و|�b1���P��q�R"��5��f�	���g����ߎN���]��x!��@"j�ݫ3Ꮵ�!��mG�nd��
��WFPƙL_�a���3��I�w��)����G���r�]f�eь"�dBK� "Q�TX/�Zr���\���7a��6ݛ=��>"�ϔ|��jh�jA@�>+�0jHl�����=� �j`֫��DW�K�N
y���J�& KP�0�"��dh��"W�+0��$�K1�b$����4�L���)9�T��Px]�p��c�+~[�H^?6�mӕg�HCqq˿n��gt+��"�Kf^Ne��$�C��7�I$V,h�����@G1yb��`���jD�
�U;�����V	�^J4}(���FRCMZ=���ץ�&���<G�J"!Q�T\�����`�. &	��Y�I;F!�Ⰹ��ڡ�����df��P��,�C�	ＩYG�쏢C��p/h%0|�{��&hN���k���`�E��L�j��⳩�Ϊ*� �QQuz�+��RǺc]g�s�*�,��@F�" �ѱ�ِ\i&s��=M�U�]��uAJ� t"@�T�pU}V�ƃY%�CiV(&�R�eV�MJkdI�@�Ͱ)�pX�c�T�VS����3����߫~��G��Ԇj����gU�����g��z�?5�L]D6�"k!�$I �Q���S�#W����J��bQ�
T�C(��x����+�:���Cjl��G#C���Sj��d������>�����SF���L���hv�╍4�����Ⱦ����/�+X�3�iT�p;��N37��������Z�vʡ��"���y�����t�~�T �Gq�AP>w������AM��)
o��9+���"�ۄ�z���V:?��0���T�Hv]�!,&��z���w^���o���x��� l 7���U0������=��f5�����7����o��]�$3C[CQ�ɐkGm��+۶��_�f�d���T@�9��?��~/h������5�p��6� ���� r�� ��������XD�Y�j1�M�;�ؼ&�&pSl��:>��y���|O�|-O/���;�]��n�O��]��	v�C�����.D��D��N�����v�MGBx��R����@��e D�I�	XAd�JI�BkHHI&`�	�[��C11���(UR�ȕj�X�,ZUZʨ������
 ,YZԨ5��V"*�PQF$�J�`��q��� r�K�����Z���$���yߥ��Zn�ܪ�݁C����;���Y_   ")�_��}]����,���xh�|����������}2*�W1i4�4�P;Gh3��G?r�]0I��U跾{�oqܻ�)�dX�;�8�5P.o�zɶF�����14�y<(�n?���W7�5 4�d�;�<�L��/1���0��
�O��|W��V}�s#�_��q�����w��$��|�u%�����}�SB�!1�SF��`6U�[T�Q=��8t}g���t��Q�L����z^;�������f�V;����h)�:O���ݮ�q�g�Z��*o ��}��0?c^�.�����C�h���o}��n� �P5	(>�����M��'�?]9�4|�%��B6>�M�����y9���Ӝ�k}�hoP��O��Ȍ~g�|$�U>��~�?�N���]�o�*� ���ʩ�L養s��������=C��U��>@l���ʱ+�����w5�~v��������{�o���[L|�[p�LU�v�[��YzN7��{�f�n�Q�*l��݇M�J���{��/�}7U���x/��n�C]���= o&>) x�A����s�g�O���XWd����P���O�=`Ep�B%�<<{�Ñ��3������\��a��'�sh!}'��=�����y���f�~�S7g�6ʛԍ����x�ː<�^�?#�v�w�iio=f��HN�0�`~�3�ȋ7��H�����4�~o����za��Jh(S���֣��O����x˰�����.�׽��L�؆�0��yM�����t��7���r�}è�}���~���6vpe�~�r����9��k��S�3#�n}����S��ޣ�f<PGǟ��k�J��nh+�^g$|�����^k�igD7"P�D"xǬ��+ˇ�!�=z��nX]h�)h!J_U�t��9�G}����6���t�����v�
�\��/w����к���mM�L'�NG��s/1�ؿO1�걱4�{�G�����=��>����?�����A���AT&�M�?'���P�� �"��):y �ıSMQBSTWd�*U`��	Z�U��B����#YYZ����ڂ�B�b �Ԩ����DcXŊ�2+�a �m��P���T�e-�ZX�T*��DTT��-*�Z���jU�@�JR514���S@�R��@R�D44( U+EIIED�QICUP�M,M	-TR�*�X1�������ɱ��������kZV�&4E�mvZ���c�a]���[K)l���Y���W��h�y�K�g���iT�����5���O�<Zs���T��%���+����qTE�M+Rڌ�eO~�GJ����q[���u���p�6pe-��ٮL��`��jĥ�����u��,��|��ZsֺZ]�gwYʝ-��m5�u��c�δmQJ�z�����U^r��mQ��M�$�	i1MA�1MAC�`����u��	�%eHW�X����*]eTY��S)14�&Q�T��!��B�kR1���X�YX,T\�HN�D���Yޠ��-iYm�����b�Q��,TTEPbKTR�FZ�X�E�Xb���E�l��4ͳm։bl��'���������(�AB�R�m�F�Vҥ2�ڠ�h���Um��5��mQmZ���5�"�U��E�+X4��X��*U(ŋR�mR�
��@ dȤ���H�(Tm
$bZ�U�Y+F
�`�T+ ��-e`�KQ-��!��sm-j�dehփhU(�DA��5(�U��mEbʕb,��-J�Q�Qj*��%�
ڤ����AQ�e�V(,kb##j*�J�1E"�QAAbD�V��EUAT*Ң+F�(ĭ�l�"����mE�[1b�II�ň1 9�\�M��׸�d m\��߭��'���*�h*Ơ'�lP�Y$?�O�P��V��-qs���c,�͔c+�:_��g�������md�V0�d���tÎծ�Q�R#�u�h�͖�S\��s���Em2o�m��j<��ܥ��%���W�[�W�P�
2҈�Y�Q�4n;SQ�h��\�DPE:�%֥�iJ(��[ݷ6�
�&��fpب�-V�[m�����)�F[/�#�W	~�X*�J)o�/���u��o(ԬhlTKJ1�m�JT��ѭ9l�ڗ6	[K��j~;R�m֣�J
j�O�t���F�Q�b"�1,PP��hn��) B����2���6�DF(��cU�Q-*�խ�%"�pQ��y�(qW-���u��	�XI	 ���!h�����KR�*����Vұ�((�?�F��AH- T2;��zWy<�~�)ޝ��������b��`��Z��ҫiQ-*�mi`6�(��e���jW��F�Ϲ���I�F��0v0bK}~�k��i�k��2��PE�2ζ=���e�����?!���+-��O��=�{�������P�~Y@�D!�Ǳ/���� �	W39�-������S[�(~��30�~�n�������_w?5�|�ن ��bdxG�?�>F ���Ok?{c7X/^s��T�Xd]�0.A����0���S��BȂm�4�B�g��6'�)��"���È4@���0��MDS"��1���33 -P
"ik8 �'E)S�*���V�T'������K!�����~߽"����_��0b�<���7�`����~$?�,9=�??��G��??^g��!\��?\R0���������&a/���PN�sd"ds1!�0�2?H~��k��Y?t�:��??��'���T('���������9�¤�7��?�߸����`TT��`~$>���U
����;�C+��9�����6�>7i��)���������/~̯����'�z��?��?:r��&��i�<�"��2~�?�O� �g���~+�ߤ��<�����+?t������ày�UW��ClYI��礢o+'눿�?��~~��}��?~�ч�����g"���C@�Sp�,�f~~�,�C�t "�y'�{��ɧ����$�2{xg�O������L ��q8���)�[)��j���$a�"s �F�
L9T��O������??��x����?��).i�$��
���b�X�����i������jT�x���~���q�Y�1��?v4���k�~'vl1?7�����q�� ̰`Mܒ<7p�	�7#��CԱ�)l����/����B�"S�J3��o���z��xxN��O̈́�H�@��/��A��^��S�O��0�p����ST�v��8�ύ��ļU1Hw@K�
7B�Fq����i��믵�������<�qI�
#���������K�<�:��y����Kg������K�$��j�?���I�'��~ߧ��C�������[��D�Oه���>%#)�H�^n�p��	�T���dO�!3P����3���7�(���������q��=�_��<��B��H���?�[�0̎�rmm-��V�jk���+n�8�)n҈�a�#Z�PFZ4��O�yЪ��r�W��5o�������d���Қ�Ǥ�~�i�N�*��긢NG�.�E�B��pq~�Ф�B'�@���dR"*�[�é�QT$A�����Mq�D:��~N9�;߬~��u�jT������cS�K1A-��9����׼[�(�����n�P>����&?���_? |Sb���"YԨ�u�(�c��S�1�k*��SS`.p��(O<�2���bȒ�@C��?�8���fH� �̙8���H�$ක��Z]ر���G��P`�i��S�SOj|ß���1)h�ҕ��>����()ey+@�>Lw��;O�s����?!Y����2
Eb��~R�`�c���P�Ყ��(wS���ߘ�l�I�ӯ�?� s�3�nS��4��8qB�nxRz��gH7�0BC��� ��	��:�
��o^ӿoB���J�9�>�EZ�vtPT�E)���-��1Y`11D4��i�{�ĨnJ�&�8Dt�bc���a#�+a�`��~�M�ܨ�蛺�$���R������٢z�RB����?�D'��%-�Z�Z�U*5h�m�i[--���c[Z��icV��w�������8��Q
� ER)++eb��U*X��S��bw8D�-G���!t����I�������@��3!P��H���2��#�_a���g�!���I(���"��� � tu>����;���ƈh^q% И�AB5B�B�"P�ѱ�lmf��˸8p����2ь��8�lX��\�.QCV���52&  6����Y�H~�aCFQEED�TE�p�O)���	��H�M"R!14R�bLKUB��H��8��QF!���8�!PC�6�?�VK=k��O���a�>���;��'�`gpn��|��x>G6��`ӆ	������J��Ji��
ZB* �������� ���nk���� q��m��%��}O_ϟ�I�Bj�l�w�]��G9�4"�iR���1VѰګ�hس��c��/�G���X������S2x���(0��x����~���q�zz=��8����Uê��O\���of��782 ����̀נlv&�C���a�A4��v��w�P���[������^���?�\dMr��^�%��.������'ѳ�#�����_��~,��4:kǇkpu�R~,)��k	�#!*�@����G�"�=���z?�����������r^K�v�$Ф�/����90��g�0$�' k'��9��]��j!�޼O���?���>r]�Y3��J�V��7���o:7����`+������& �����;��?����N�Ȅ"8�22=�+~�'Nv�6o��3�im������~�x������=C��?������)�Y~�?hߧ�Å���C�go�d�d�_�?���I`�9�C��#�����B�&�QVq�T�0e�����E�~+�jSq����gᎏ�>u���'�
���阣�]�碲��l��ת~�������{���}�s��&4+���6��ΨqBT� Ed0���T�ih�kl1�OO�p���sH�R%(��4�lv����l�!֛#K'+ak�c�����`�0¦	$��`O�NH_���*H~����o�B����ǯ��wb���o�m�ʴDƆX�I�R?�a�D�h�f@�7��\7�h�̘:C�A�c\Emw-��gic�mOۥv<��K}��@~��w!����xg���L��C��{K��.W���0��ɶ̟K~0��0��PZ]Wy"����2ki�	�|��6 �	_sQ�r��Xۤ�$Y�K8]Č�#x�;RrC�� I6W�㷽4�Gƶ:h�#��Y1�x����_"ҏ:P����l�`��,��m�^�kv>���� �@'�/���ׄ��Ǎ�8.'�.��}�Wgd*m�]����t� �( ~�Ⱦ[O�3���m��7�Y-}����/��T@���G��?�8�c�����o�O����/���M=�Z�֓����}���dV��������?o$�`Uց��/~a��,Y��RO���EhG�����:\ݫ?�8���ﱭ��R�r�o��sy:Y����뻾�;&���S�H�*m�=��T}T�K'�\�e��Le����5�<���/��?�xo�=.��>O���!�~����~UPy.� ��6gK��s�������x�su��]�����_���p����2�b���N� ��!��R�j�:}�;���k�~��3��\I��.7�{����>������j�Q�O@?w���󼧃𠏭�C1�#��������������c���''���Ӣ���.��� �L}_W�-����g�}�nf���Ϩ[�2��p�V���z0���� !����|��hW
|k�s�`=4��O��>��\�9������k�� }���|���V`��J����[����O��hf]�
	�u��s��v��������!��y9!.�T=n�_%>� 9W�偰@�'��7��M����--�}�	�M�q�v��ᨩ�@!B
P#O������|��|4��$FP	�;�20�#�bj6�o���a�~�j���c�c�{l_ë}���M~Z��z�@���r��+�Gu���` 5��EN����јu�?�y�ى�75����p{e��sQ�! ��k��dt�K�1��,���N��v��p<ֿ,f9��w+e�喻S>��A�c��q����)�v����ݽ!���-e<����*�@E(���*���^�"��'\ڛ?Tsnd�|�X�C�=��9M�I����E�㐑������g����vIKЎ	�	��}Ym���ާ#��4��Mτ�b*�񢈭#8�;�d�O�~�9#���K�e��2���>�s��>�֙������^!W��0�}�_���m�����@B]��~t�]�X$�12J_���M"�0#�$;ǣ l;�Z���3�{ޞ��������ѻ1��_���x��7+�"*��a[��N�f�i"�!;Q��J����S�~Mr*�������a�Dd.O�St��ؐ�6^3����k�#�Γ�a%(X��?����U�v�?&���QPP�ΣD�>��J����)r)�*��2>�M�'���	�1��hbG�^�������O�EUYsɾ����C$����I�ڕs�Y'Ǉ��g�:��t�Va6��{_���I������~���o����]<v���7����]>�[G��<�=��O�:?(�U�:T�����y�{�O�>�\4��>�B�:�zM5�/�H���Խ3�X�׸w˷�(0v���Ў�-@���$��[� ���W͔:���w��ry������ h �ڵ�A�'{M�a�d��]��~'�}GS�x���1�m���������v�����/}���|�~w]�]�ňp����qJ$z�}�pp>,=R������#�p��	+ьG�f_���7z���P��/�%����g+0��}�`��g�!��Ѯ����j y6���2O(�ι��^}��Ӽ$v����G�p�5��'����_��8�J�!�IӬ��Ż��ڔ5�V�n'1g1ٴo��>�:�Ca�|�l�����\f����~}ӹ�����$Gr ;�
���E~����HO7'���{���]������.߷�����_��o��������Z����r������Hs�(��6O����'��������bR���|!Vr�f��&�n���u���:��7��ؾ�+�].�#�߸���������Gmvk:�~H�W֑M�9�8?ۧ�fq*������
��a?�_�����՟{k��H���*�؁���]\���}m�f�=5:�\ 2�l<�yq����:�S�þ�<jcMs�؟Z��'�=���N(G��- ��SI}LȦ��-��ۚ<�*���f�Uܮ�����rh�F�pU)K{ѯ�*+���$W�d�"}:o�"��&1��pE���x�";�������M���̘ى�&[Ճx�WdVe6���T�`o��S4@�9j�o��/
�7r��.q����ۍ��ɂ�s ��3��'6�6��]t[���f]w��߯���w���!R�r�]�3��ߑW�d�G۞�`p�}I���/�N|rGM���?%��4+�JRHZXB%Q�Z�
@�{��(%�^��_��(cH�.�z�
�>s��g���@��~.7fNc��ynO51�̗Q���vRJa����!�ݎ3�����s���7�CS�0��\��I�h�Ɲ���X�u�����!*��"R�("`j*�R(�j(��*"d��ٛ6�`L�V��)}Y��LSP��Utz���Np㌣A��5J����J���EQ��=���UJ�+mUZ0b�l�h�z՜�*��ĭ�5,UQ~~�F��x��Qت�K�~��U�ܥFڦ�U�m)l�qr��E����^���*D�="g]Q1�QAQ4�4SQ�PXG ��?��y\�:�ٍ�Mt�N"�_H�];��.҈\5UPQSK�ETI3D�LTRT��z>ǱBt	:��US*�FP�*p�mw*�H�KPjĴw���Ix����Z���_��'�~�9PD(��� >J	e��à��(u?�E9�f��������-)p���Bm�Z�2�Q⿟wێ�;���ڣ�w���mu
&vhV�wum��Yv�6͊ݺ�zg����%xS��G%Ҍ�W�����Rx�Ex��C���u�ѶY�H�B��(�����k.q��U]O8NN�����ˏ����W�;)ڱ�+���@	H�w"�:�r�����e6�����{���`ΚXʲ�2�j�]�EKiu��]��fښ�q˓��R;yJ^��K������ۢ� ���K��x�${I{�>��#��O���?`���wI��7�����
��/��*�)Ꮝ���D�s#����Z{ڂ��=I
��O/A��8���T�ܥ����xur�>,�;V'��=O:��s;]>���%ҽ�^��.��fl��%4%JҔ�@U�a=GNș�U_��q.C���6K_�z�vU/�w�\W�[ ���14�Ds���y�4���&(����
?������"LM30SISS$�!A��*�F�(ƨ* ��*�X�(j"�������")�	ۨ�{�P����p_���탠<�����F����:��c���e�O�h���>���@�H!�4�2����0����T�2�S�R��W�*w
�:��iU#�;̓�q��	��G��N};�0Xz3a�i~���������10D������1E�9 W�\�8�P�A��G5W�y\�G2YU��ieW�龓�\�s=W�Ju�7=��WRr�w�/�]G�;�Ҫ=L��i�x:�i��p=��H�ƒ[Ux�Sr��<ߔ��s_#��D8���p-�	�f�ܣ)s0*l�}E��d̙��a3�jn|F��𧇫���s嫸�Ju�~m�%D���b�ʇ���g~�+�����_M�)|Q^g��������;�ᓪ�2~���aU�=Z����yS����͞7��A�xk�����*��|y�:Jw#�T�5��y��/��ޓ�;�� �И%*�� 3S�4Pr`��5^
�lf�B�>����{u���z���	�I!�̼�����W�=J��G��gt]�j��2�u���9OJ�ʮ�>�Q]w��2m��!Pxj���zO���Ooi�?�7����u��s���)@��`Am�X-j��E8d?����Gi<ǻ�jj*mƀ����B )(�h�TP�O�r1��߉G� O���"H�����)imQ����VMc
h��,��0�E����m���:�;Ĭ����*��OZ�`�cL�z�0�6q�5: ��+��|����f�l�;�c�)}*r���;��FE�(�8%�M�V1�ĕ��q�P&8�"B�T�Ь��U �U�mQ��kV*�ڌUY`��UJ��H)Y**��F*�YZ���F�"�� �5CT�QQ"D�2(�(��UPJR�iD��
V�*��El!A��DX*H�i�b��(���f*��"��)�hi]0N��O��|N��u:��x��6�k*��H�) ��0���K������W�<�����C"<J��}�Q"�%�?pG��c#���6��*	]�B�}b�T�J����G��S�ҝ*�������5�>�W����}"xjrx#�x�ݍ�����T#�G�@��o�N�s�;�{A=gh��O��S�����	�<^Y��JZ��h@/���g�����1h�i�?B��<��/�+���� ��B��3��\��&64��0H��\���{�i����7�w$zY�s��3~�	�|�6?��Oo�r��}^��~q" Όo��~���>���O�}������e�����o�]���� {W�ܔ�;Ǭ����p�h��كs�Wo�:`��@�m  �����<������O��+�����P�Q�"~��̃�;�{��b�q��W�n�.���ْ������ޒN���pD����6S�M���{��P������J���d B�1���K
�.,��Gx�S��˗�:Az����꛺x���,���wⷅܱ����>����������#_���M�2��G׾�D���pd��|��`�����8�����g����<���^�8�XA�/�v��ga�ҹf~��m-c3�3�h�?A홢��g�)�ĵd�Y}s�<�)1�����༠
؎EȮg"��0�� *�<1�G���G����=?���U���_>���ETC�#d���_��~�~��e�cT���~�������N���G+���Vj@K�Z[EP�P��0BK4���� ��1A\e/�`lo�o���Ib�k������/�3G��6�sy�O\f��w�Úm�ݵh��:eYY��]�O	��������G��H�P�;q?��\ �� �{��O���PG��>�S��K�lw/E��^�_�Û�j�#�%DDO��X��1TK[HD� k#��jE����<��neV]����J���U}F��+�vW�H}J�d�˧}~��:�vP��5Nڂ�|)�:'8�	s��pv�w��j�M2�\��ت���UvG�ڟ]���<?'�8v�?�o���S�}>K7�����,o�����A�K֓�S�������	./��?�~�E�~pa����ģo[�X��O��Q!�?�+��>��0[������%@���͞�-x
�H
���	=�{�X�ޅh��3���%G�O��d��h]��ح�����Jb�����@1�E�.2�EǛ� �Vp�&
�
�P� �*������<�2�D방�͛���FA�+��������b���������o_�z?��;���vc����c�w��?���w����g��������T�$z����F+�n>�>��z����zs���
іߪ/�Ʒ�~�����z�_rO	����_kד��������o`�27	R�����g�}^9�}ݽ�/��.��;��!�_M�l7������ⱃ�l!��b��D��T���x�x��4��!'��K��g�4��3m���#��.h��G�U�m�-}�{Ǳ"�֯��[��� � ���f
�&����*"�*��CF(�b���IR~Hb�q��[��|4��5-3�?8O�Th�O�M�
bW$u }?��.��4�����kw�����#r�Dq8�7��;X�)��-�a���9�mim�
�)�VX�c0F���G�����~?�s�{���3��5��<׫����c�F���z]����~���6�KKe�3�cτ�o�II1E554L�R\1��o�o�*��PTHQ��R�%)AE1%45�HU4P4�p �*����Ӯ�N�U]���F�#��N�O5;��j��A�KK��^b%�9�����\�}
��Tt��r�:�9�#qC�L�	^:��l��hl��NA����]rH��Ud�_v�8�^��Ep��5e;��]|�{�r��A��|r&�8>����{���4�������J�~���O��䳯�e(�w��WӜ�
���?�+��?N��!�U� y����eEx��NeS�^�TiN*;$�����*8�n�E˾�z��?��]u<}�o..�r�j	�*�^�s0?��@x?���?��3�	�.?���$�1�ˏ�19
��UE��Q�k��c��pb��`�E8��(L+Zj��aq��q��~�N�����M�8ij�hi����f�()B"�iFA�E�TW�Niqu�/�U��n�u~B��R�k�=�݇�}��*�t����=�����}w��hΔ��o�$���:�@�\�~x�}G�/�U����5W�������u���>�!O��[����|B"�l����,���d}>�Q�r%˚u��iaHffC�%�I��M���Q�ph�JV�f�1`���Ӑ�
|�B�SԦ᭺0��Q��� E,d����pX�m�}Ӷ�]k�M�r�����"�)�*��q������?�Ȧ��l3��װ~�)�8�SE�UUHDQE����"56QAT���;�=��D돢G2�'/�}}�9V�:*p�_m�)�k�p�Y�(��g���J��t'z��:�w�<�N���>����/�4�u��s?s��TwV%��jBG#�yxxty9���]�)��\�ǎG�p�;W9%�v��~;��W�������2|�����൴��MU4la��o���b��k�Y?��KI��VS*Q��M!��]칇�K٧(���M\�#Ӯi�S�����?_���}�G[ڿF��K�I������:��I$�� ����������91]�$��\�K!�8�8bH��.TDI��o)e+m���?;�}��ˬWs�l�TW��0������wsqt�c,dcX�1�C�����}���/;��_��>B���/��>/��I�_8��p���ϭ�wK'�!��0<?��}�)��'�(�����CUu�D4�_��rB�d�� �9�n��@�ӌ�gT�K�U>p�7�'=]Pi9/���-�l�Z5�U�N5vr��c�:����>���W[��-t%����~�����9UG��Jj�[���^�U	*�U����_��w_o�s0�������^�ȽH��I|�_����R8%�?}?��=7t���%}�OQU�]�N.������^���N���'q�\�l�(ڬ�Ey�6" ��ѱ�p���x�n�o��/z߅tò��lqO�_п6rs%�{���Q�yn�9x����t�V����&�!�{^�=��2���/c'�UHʫ������ȧR*�������/o��P}�5�֯�љ�:�Ee$���0 � P��� ��|�Hz�/�	�^�X��=��)�$f�!��^����]x�h��e1��S�]6�*⃡��@����~W�As�Ļ�.Z<T'���2x����[ ��{���us�{���u'S�M��~���O��w�FF���:N���}	x\fG���뾬�L�-���n��p�4����\�+���[�/�S_�@yD��?��{��g�#��r�'���>D�M�>9ܙ�q��r%'�!�8&��p�`���"��"�[2@���0'�#:l�O�_(�����j� ! ���p?�#�wC��Y��Q`��0���]�������m�%^K6/������w���?�hf="�G�,J\���#�P�s(��VF_��������\�i_�������󝈼{.Xj�~�_��Ɍ�7�k�*G���MH�^�[�Ƕ��f����{m��\D `~��M�Y#�J�R������_����~��{^���=�����>Ϣ�*~q����L1���,�?@���}�+B�˾�'�6����I�k���� ;�K|Q�	=����ҫo�{#�*犢Uu��/1"�H���Q�%S,�B �"6�� �A+T���B͔�E�3'5wf6��O$�ӽs�[i�¿@,�2"22����E�~��W~鏃��ie��=�j��H�(�<4���SQ�f�;]XN*:�]�	��|ݲ4�$�S~�.K�}?��F��8�ȑ�����@A�@๋�� ]2���<�����������{�򿯿o���i˞�aM����4u�W�x��&�J)�/��H���%~׽qs
�qn1j���uA`f��&zO#G�u�}�T�+�`�
�i�,'�dk�-q���"i[Čcե]H��K.�+�q��]�&��	Ee[���ъa�L����P��)n�Xy�)%�p�۾Ij�:^%	�LI?��`n�Ty�/	�!zf�}s�N�1��o����9p������vG0Iɓ�r��`}?g!������h��P�'0?��v;�P�W����cQO�/��d�]z�Q@H}'q��A����ՙ���ys�n�S��t�d��3�O��O���m'L ��	M-���C���ڡ<3(�2ӈ�h����o�Z*�":���>���*ᘊb*%iP
D�
}$����~���w�>9Q���u�MTTA�6*��h�("	�����GP�?��]�0�8.?Yȡ�	�?���4��M	��[���đ��	~�c���N�z�7)5�iTi@.����C��`N�9��k����f//��S���SHOK�e��_#�L��XMN#�V"�aO�@}�K��< w���K��I�$	�ҫx�/�~�?4=��Lk���H��xטj����	��C�!���=O�k�s�L�!���٘t$<�J�#y'�������:��O|���"zI���PՄiQ�
EO���;�~�����n�;/���s��.S�|��pr]��"��9q)xI>��T76Jn>y�߰<��I,�����@c�k9��^�_��3�oP�(�G�8��!�~o���%������),��<��$=�vr_K��5Fz�������`8�;�wP\�2Շ�{G���fSְ������)QBu���b����zv ���H����L��a�@�&ՠZ ;>�ϩ���<�i�>�ޛ�yԾ���
3����W1��~����N
"�~�������\��O���^�)����ؕ����yտ�~����S��_�S%�Qe��W�w���Bf��}�fa���9H��K�w��?���	�	���ܕ�B�Z"G�[���E��;�y慄�(4/kc�3�]r��@�Bu��g�J��:DEo�Щ���\N�E	�E^�<�B�t>��}�2�H��۬��FD�F�3������翎���`Ї_��"���]dC9�WB���/:�����:�)���_3�LUѮ��a;r��Tl��5�X�#9���rY��.�$;��gB�֡�/���=����jυ
�3��2h��=vnή#������7ܝ���9�
o�� NjB�a���2P<Ԑ�VBy �f~V@��B�TR���b�*MhF�h@��@�H��q`�^��{�d���AghZ��r�)λ�ͬcm�W�4��q���2v��M@ �{O'2A�-����+d��Қ��~��������� �;�<OA�xN���>�xO��������}���OO�3��TވE�/���D��S��dA�N�άDL�QD��Y5����#����4��z�5RHT�,���$lR(� ӈ�R1���J�~a�\s�^�D��w���J6A�T&�M5*"�׊�ŷů0��+$��BVzk,�G:#�$.��"P���C�������I���Srr�8v�.����N�������9���\���_Lb���_�nl���*z����x�����"�m�˗��|s��{x���Wh0=���IJ���oNkeH���S���"tE��2B׾0�?�j�M�/�f	DTW���I�=���s���M�f1Q�bL�F��*+.�k� �bAP~���C��/~xY���Z�m�I��`���@�D���e���音��o������������5r������э��]�ZZ^�1�w{���c�*��?w�&�����`����ﴺ+�X�z�KO����Ե|�v�_s�74�	��2�HI�$��=61N��+ ���M&z&K�T�ퟆ�Y�}��U�:�����O����:�kI��{c�&I�����"�����wL�~�N����c��*���� 6��_���z�8�?���|>��޷�������I�}�C�����*���
������)��`���N���y�k����PG����3)h �MG��|����{%�;���=���G�����;j�k���O�����w����u�����9���{O;���Ah �����闆�|�����?czSa朓H���{�wٿa9��4%O]��S%��eXM%���?2C0rAbu8t��ZD��
��z��Wu0�@��[���5F+x��Cy��-E�� F��*�
��\���c�9����̭�-5H%hO�c����������Se39��I鎨�*}�閭���d�
~P �I�=�⟑���M����#W���K1^?��Z2�3Ȅ��b�JmX���!οl�_�?d�`�H؟������ω�px���ج��B�H��r��@����q��Љ/ap@������@g�~K��\�S!��F����$�p��?Y���v�O�2�5GSM�A�u����={�`�@S��21�BCw�<y�Ml`��q_KH<a!���'ؾ�c�.z������l���>x�i���i�	����1�/�w��W������QR�d�ҹ~ ����3���=!��uR��Q>t��d6���5M��a���K�sJ��+�e=�Q��q�q�+�`6s�R�C������p0����D��A�'w���S��~����W7a:���x�eM�������_d��
�߷ x�N�!�Y��.}��u�$�\��̚��L�ta'��Dp�b��w
r`�Fԛ�(�� �L����U�~l�b N�ǌ w�����i&��O��\��35t����)�&�_�Ü�r=���X1�7zHr�%�;��Y�)���e��j�|6�>q�sbj�)�)G/i�>o��w���0v�&���������r=w�c��,X��Ogr��_º���������dy˞a��i�͸D²V�&I�6�����+�N�?�nk�,eh.LfK�}�><�>��8�,!B&�a=I�#����B���9��;��o�*�y�s'��$���%!0��� �h�b�5-,��3U���xl��9��&L�0"_�:P��NODb�C4�V�J�gW����?���^�0R]Ub&D^?Jo���B[CU��ej��j`ɑ��j��x}^Qˊ�����V�4�	a�����1��h��\C��Ka`�e��3M�݇���A���u$�5DV�"P	N����|.�>kr\�Md�`�bҵ52��22b@t�	J-+HR#9"d�Gb�1�^�}�9��WR�(F�d[�ll��T�j4I ?�����u*�T[,�D�������/i��g�IeP�O����yg�k�`�$QSD�B�0�� ���^�׏��n��y���!�U���g�2��yC��k��t��S`�2�@0�߸����	� @.��??�EwXr�jn���`�36XM��^P�J�ȣjB�1�b�m�qڎ�e��DB��LSY���2�c^�UVI�g�v?������>�pF��J�����/�,,5L�F�U�,��S ?��;��}�KE�Ӕi�o�N��`��.'^Q��_
i�B�4�Q�`�wJD�)�=/{Ibu��p.�gzY����ɣg��,� ���R��@�g���f�Z�[#"R' ��~���"�ԇ8 `V�(F9�
���{m�ϰm����;|ٷ,�4�~�|�X���97�p�z���FM��1�ʰ�_�8K9&�}u������bӼ�<��l�+����D$F��j8��3�ҧ��4wL�B�s����c���`�V�X[3|P�����:Ҩf��q�gl�6�c�͛e�d�ƞ�=�3�Uن0�@$`���,�|W��QhW~c���ѳax�W�rt><�LV���xhg�jE'�f�+���.�=�jf�}w�Q}/�Hϥt�L�i��K둮��k�}u�)�l�����aq,G6�xf�c��M�C�oq.!�M�Űә��
�l�����ڸ����c}�F=6]�!�8P [c���m8�8�@C�Pe���e�P���:�l5#Hi�i[6l�ƕ������UmU�2$M���
��+d6�Hq����%&� $(�^�m��nY�g��s�[�+8��x��<�֘����ѽ5/?�-kÇ���E��։�8�}��S�\tި�l�X��u3��\�bY	p��rm�7{�ߏKϛ?��r���Iח��s�xӪs^q�l�r�6��]eۚn�=��1���7�9�MJA��C�ˌ4����N��G�1�?n�yg;�ן>Z��x�u�(V5���l��y�*h8S��x��kY���,iJ�r�#"6��,qK.ت��G -|0�գ@ ����}��.�WY+Z��i}���9fS���D�Ȣ (�Ԕ��	SDUTDST�QSKQ+URLQUM D-	MQĔ�MY��YX5d�djb��1 d 2 `��z{w���<����C������%�򷍯���>�ʹ�'������:cXW��v���s�6ӆ�����[|��缟H�myg��N)8�2r�;.�e3i�^	�i�%A�,��t�]!�Q�W1�NP]&�@�(�L��yd�3�;e>Ps��v�#�u?�\���>�=�ՊS��8���a��u�P�kT��Ç�.���צ��9R�<x�¸�S�$���lG���b��`v�3��u��m�|n��H���y�i�^���wZ�˿	�������x����ejm7mM����� x�)�����_����Jփh �@ Aj�  ##!+�D+���	�Q�z#���YrHQ���,j�e��N:e��0�i�@!���u�Rǻh
i*��#�s���h,Z�P$/���؂�� (�	*&P-q�l��UA�q�aTL�af�z"y��PI��� ����ÞzH�e�L���Y2BOlҍ�
�b(�������6�x/�A��"`e��E�BჺiO�2�2i爲���N*���E��G-�"(�	Dh�(�K-Vp���!C%D������G��)��DwJ�t�9r彭��/.YK�X�����S\�u�]���-U� ���6�-�#b�K��q,ӊ�z�2���Oe���-�o�mwm�|����<��x��7w M���0� Ȉ��}ּ���o�۷N����(G�}c��A�J����ʊ��a���ٶ�CУ�$Zf��AD���k�y�4��Ev�#����y2\�IR%eB�x�,ҢJ�+��'�b���J�9�4�ڂ��*���E8���AY��rc<��x%%U4� �<���-�iM��fh�L�N�D��6C���1�B�S9=<��S-�S�T��`��26�E�R�!�	Z��E2G!�Fi`l��4�z3����1��)A�B�H�DrHVK1��
ꦓ�xDY^P�W8��}��9zl"�;(A9�Kq&h�R��Q��9	g@)8�4Gʬ-Nu��(��bh���-��0���gӏhZ�D���N�Di��x������_���~g�g�Y��\�����`��U\91lUBR礨�\�>�`	H�t���n�p;U�Źp��PKq40�AaD��da݂#�h�n�]��r���Ȣ���� �a��j�aPƌ�j�q��PI��1dd�ClY�J�"eB�!g�M$���S㬴G@$O?T"$��z�+)���=]%#^Z�}���Fr]D�-�ۃ ��$�/��?�Y�H�
)��AezA\��Yp�� � [�������x��K$�
�2��)�1c�X��bU��(���PX� Ké2㲼$ȍ-�/���%[H�]ͅ�Ă(	"�Hde���)�HP*7t�A�1]��F�q�B����-�IP��U�	LF}K*V��H�y-�(�L��q�0�nL�_v�ݎ`�3���?��S~$aR9SE���hj4�d���1hb���a�SQ�� ��i�$�[U� @|����KD�g�!�>G�%��)%����3�7.��QSXԚvH��"H�4K/	(ŗcL�y��T#&)�u��K�!�)¸E��f�NZ�Y�`iS�����L6ʄ�|�W��	\��}$OJ!�,�]2�
�5eDGɦؓR�&����B�����r2��dN���C9D�8@Њ�R�/Sd��q[�y��X�g��_�Qc�d��i,t���Y�Q�� Ufhu�˺H��Վ��K}��:l^0���\�ՕvFW)�M>���l`Ca,���,''��z��͗�57y�
:���5	��XYer�QK���C܁&��"t�	������-��!��#䂉�<�\}�V���5��%JNJ���vP��d�9��RZ�H�`'	4�.���H�k�ɈzE�>�d)�*	2	��o�����~�l�����i�_/����������z_,ߘ����{ߡ�Y������|΃�9婎�������/��}�t��l������֤�'��~�+�;�~�������{���I���Af����u�-���Xo�����D��.p��8i/_�>6?�� �a!7�?��e�wa�rc�{�W$WH�&����~����|U��.jE�_�����\�������^���s�����=�ZF�O��s����n���'t!�^x��О�����`	�p:�{���z��e�5�&ϷH~�wV9�P���;A ��P��{6� �w}��)Dn���D�&�rR'R�$1�����0���ݷ23"�Վ���Z.��\C��V�U��Kwc
�ɵC��=�J��o�v�AuG�jZs�%F��QIK��c8��\�oNee���Y`pΈ��t@�ʖ��҅�@QC6fPEL!,�]�6��@�~aH�\hlUو��+U/�-­��m�,)�CJ�a�~���;v5LmD��� �5�E*��	� ���QTA���8���(᭕���t��$i�v�(�B�����
��C9���U�V-v�ɖ}�s^�5E��6� ^�5���#ްɉb��L�1$n��[|��*�a���Cr�� ���� �X�&
��e1N�:eR1�aa�y��60[4��Z��������	-G0~("�]V�B�*=r�ӤP��~��-M}�-�C��-��ɯ(,d�y��.��Wm�f�r�x�L���^�����3��UP�@��@ Z�h!�j�-^nrd��ُۂ�%f4�βhQ8p%�T�d���JT`�����UA�a��f�zf����O=hFm��,�(��$�Ҁ�#���c�9r츽i2���=W��5^#K�Ȏ����(��<����Ӽ� ��6U$�,��#w���1���Ƀ�1$r�Bv忔C`@XҾ�"����e+��Sg��S�XkU�4�G��%0"p�!���P��	e��:�v�7��RpX�F��'�0��O20��B�#D��d-X��2ڪ���y���!�[�����bqK�ǁ!�Uu��YB�Cɫ0��,Yͦ���~D	�[���f$�q:s�Yc�S3xdҘEl��z�X�	�[�P.�*�%���*j��.HJ�I*�q���,��+���c����Le�C��`���k��6+��m�@^���,�.r�q��'��e����i��D���r��r�R+���L��$���j�؃�̕x���,���3^��K&�r�p$��]�ܼぐd)ˈy�?&& ��N�6��mw�NW��v���L⧷��T|���>�&P��� �
���'��I��#2d���p��Y,Ŋ�R�8�Īb�8�L�����Jm*Vң8��$h�$�$��N��m`擖�i�mZ��RŅJ# �
��T�� � �))"Ui�W)8�[%�!�S��Ɨ%-�6��0.2�̦e�4T�0\hmK`�C�m6�M�ړj�b3DT�F�ٴ3T8���8�?���[6VŰ�M�l�&�KjT��)KX�O�����G(1�	���R�r�ظ�<S�mS�Ca�rC?�!��
B�X
B�3@�YZY�*�U%#*���0�B�*�E P�$��`V f4�*E
Ʒ2��U�R4�ݦkc�QFӰQYm]m��8�?���'���S�=|��AcFZ�q3V�"4��í<T�gjU�������c�#�x�225B���TUHR�LE(�E!(PX�%�E��3%E$��Z�E��IsND3% ��%*
AdY9�AL�m�R(�R��4�T1�RR��QD��S�b�(��ŔdJ�-R�L��Y%aF*�E��E���!i*����)H�J�j�
J
�������"�*��ZF���(�H��T�JP`�qQR�QI@U)IJP%4D��AE)I�S4PR���4cV�J(
R&��1R4�b�Ȅ� !��3����o�������w��;���m}G��O����~��x}W�����_�?��k�Ӷ������w��kGz����ο����X9/U����帟��)t}'�?��~�'IG���Ǉ��������������-���?��X����/�����>Q�o-�[�>��Gޥ�/�����������Z?����y�'���_ĩ�y��կ0�r�&!��7,��(��&Q�b(*"�"X���hj���J��
(h�(h��bJJ�"���)(`��*Z
�R���U"V	Q"�hhF���J�R���M��PڶShڥ�"�*���ҋJ,��@ĥ �P4IM��e�6l��-�cj6�kQ���Ҡ
1Q3M5D R�L�l��.�h��ʖr�d��JJ���)�cch�[M���l�hE�� iJhh(A�
R���V�)�
�mЍ����lU[U%�)�m�6��l���$["6���[�mUm([
l��Kj�؃i�F�l-��m&ͣe��V��(���h�>� L�h
%*�JH�`��"��U�Ԑ�$PU��!������j������(���j��"�����j������)"��)�����Z
���[p6��i�6�m%l���Rm#e-�[BڣiM��Ѵ3#j��������iP�E�V�B��h��T-�l�m6�6���eCaV�ԫb�m�ɰ��
ٳ2��e��f��8�q��'K}¿_H7"���r1���"j�IrT�� �� � �<���������Y�|�0O��b��[��t����^�۟��}�i�����3����?����C�����y~���C[z��Y�y��(}x�/�v�Ӄ��2���x.���$O��>c�q݇���?+_?�y�dw��<���\ ��������|���}���R~k����|��?g{�pMv_�����{�DN����V�ϵ�x5���7���v�����pts��V{u�����q�g��x�o����ߙ�������Ø�9?��>\�S�������n���u����x.���/��,������v�����.v]��u�g���'���n�ǫ�U�����Y����{�����,����'�����6��y��������O��/�]�{�L�{�)���ϳ�����|?��=�A�?�����g�|�>�~���?�����l���|�7��W��lg�?7��<_�0%_, �����2��Z|�K��s��f e*)�)�(�(*Fbe" �jj� �"(&"���������bj�"�"����"*i�j�bf������*J)h�����f ��*"�%���)�*��&�B��*I�����"�b����������&�����
jb`����(�
� ��j���
���(��� "�*���
��"������h�*���I**����I�*"" ��"I��j�i���h�����&��������*jj���h����j)����)"���*��������H*������"�����"������&��*����
���J
j`*�h����((���������"�""���%���$��
*�����i����
d��
)�j����j*)���i�(���"�"���(�"�)�"��"��)���)������&�&��QUPETQEQ*��h��)��������)�������"��J�����h(������Z����&"bI��*(�
Y���H"$���������("�*��
�B(��&fj����&�"(�f�	�����������b( ���j��
��(��`&�"��j*"(����(�����&����f	�i���J����j�(��"(�*J "J�$�(��"��*��*��*b*	��i����`�h��*j((��(���H*�����(&�*��*�$���b���� �*����������H���d�*I��b�h��I���f"��"�(��(����&*�f� ���"(��&��)����*��bJ�� ��
���**���&�"J�
� �""�*
���(� �&���"Z����H�*b��(��"�j*"��j) �����&��������*�� �*������&�������&���&����&��
�!�����j"*��"��*)&)���"�jh�&��)���(&***�)j��H�h�
��� ����&����(�F�$�*�����)���""��b��!�(�����d�h�-�����ԋ��[����k��]gu�1��E�NӒ�����������?���;�K��ǚ�Z����������|�s��s������>�������s�vQ�Γ��'�?i�O�uoo��=	���_�����W�jU�/7�\Tԏp;�b��{gII s���~�M�������oG�?����/+�s[��ط���?'�����]ז�^�w��~���xټ�?#�)̘�o�����~���?��~�h�_�۷�?���~>����}��U�v����y���M�~�����z�3�����|�W俷�/����?�?���σ�?'���}�s���?wĤ�����\�CG�繿~wg��g�'���F��� Aj�-��~�G��NKI辘��_�8�y��#���/���ƨ����al�������B��ߧ���z��o��Nj��0r�O�|Z����}JӘ�2�	WxJ�� '5%�(��U�����x�>c�q/�;:�@!f�� y]VՒ0��J/��R�c���Wt��0��
*s�B�iΥ؇���S�XÊ��� d%�G�6T+�-���y�4{>r�e�uNI�G̐]Ա��E8hh�'P�y� �˦�zr�UAr�!��3Ѐ�LX쥤.����<�9�;��h��i���B�9Y��\�ތ5���N]`ңͤ�k��N�� `m@�S�ۉ0��Ac��cL��,��G�� 5T>97��U��vC�(�jF����e��\�"GCC6�Ӏ��V�|S1����r [9n[�*����3\�Sp�p8K���	�mW�<V��o$ t�1��4�H �LY�A�IP��OQfO�c�8=^,[n̺e@i.`��DΉ�_=�B[�م�����,���O�U�hԉ̂��t�����@������7���7,���-�D�[%��XZ.�*2�-�Rp��T<�(� 꺀�&�J�N!�i�+/�@�i;#�ξ�w�ǖc�Wv,&�K�[d�5,K���,�ιuv2�şIk�U/�� ���:�����i�\�j&"�sC�K�p�{��r��,|}I����%d�,�_�>s��տ���!�~$9=����|��<���@��̓���O�<���v�����˻���>H|��� �3C�H~'�I�ޤ9����<���0>a>a���C�$����J�ԕ�s�0&�������@�'��Nk!�B��a��C���٤5rByO~�<��>@9�<�~��	޷�k>I?=�k!�'��^d�j|�����/��~�ā����!�{$��k���!�}l!9��DA�fR~ �@ "�(�mI�)��ju��C� _��B~v��!� |�W��$��߯^�՟2�Haq˷�]����vq��!�u�;���&H�3�	��;Qa�>d$���?o�'	�~��d?I�(��!>O��쐞C��� ?��a��?vK߶���>O{bW����c��?-����O�I�~a�C9���Cח����9��?�>���~�2N��|����B@�`�\��h��4�TDҋJ[[��ʶ�mD3(�DڛR�z�Ъ�ʒ��J�����R�A-�B["��٩�4�U,�7��T��s���*x�C������!?��VE9_�2I����viS�H&}�!�T4�3�tʝz�.x髦S�M�z��d5�o���C�ɘJ��$�
�瓦��+�F��nN��'��0�Շ�@��(y�}C�;�I<��0�9?fJ�'�s }"i@g�ՐӁt�aJV�D!�R�1�&����.!kR0a��� X����r6�@�0�2f~��\���Ƞf0�'��@X ,2y޲@�0�~0"�'�?d�̬�Hy�	<�~���
Na��-���H�
��FR�$1�&�d�5'�Kh6٠O�����)��Y�ا?�����������������������������������_� �[�v}�c!lZĒ7]ͱ  �P���(�8��cPE  � @ z��          �           P    � h                 P  uL    n��P�(�U OF�U$Pqi�            Z4ޔ c����65� �zn��G    �`hP  i%+�P(���{!��@$J	)E�([dH�BF� �    Q�  �g�    @ ��� �   ;  3�`    �Rg|  l     �*)[��   6     � 7���    
��<                                                 �     �q�     p�cр���p�|]�$EP ��@
    ((R��"
(D�������$R�@��    �@( H@ "H�� D$��P1�  P   @U�V��hk -U,Ӣq�h�e��u�CP� �v�  ��^���   @  (    ;��$5 ��� �Y�   ��h �@�L � �b��`(�  H@  �   �� q�P@TQ      &�  ��S�v�>� ��       ��@ a20&&L��CD�i���h�m@р�h�MOBy0i4ɩ��҃S�  �	�MT�O	���2jOORf#�z��4���=�h����OP���=G�������OH4�4zM�a j��(B�)�SM4 H�h ����  � h                <�)DI��=M=@    z�     d4                ��I	&e�F��4��2 h�� z�    �C@Ѡ    h�    4  �HBɠ ����4d 0� h �`F##ѓLM240F�0I�d�&��2�LL�&#!?���˰�䨎�Q�6��;V����Hy�u��c���0���͛B0�]n4"�����7w;oi89���<��M��N%�ée!�zғ�ٵ��sd�FF�,�L��6n��2��:hn^2����(n��O[�	У��ݒ��4���f��坛�8�3��.���i��&��t�Х���Xʶ�b�>M��]3M�vV�:e�Hm��x����Wg�\�M�S�-�pڈ�[p	8b���5�����x��Yn0��5ݞ��
�1�*l��T�uT�
�i�\���8�ۖQi'�qt�q��:b�N������i�A�Ck�"��M���_�5�;�u��������-�vx{b�����4�h�������^I�e�1�ʳ-���	�=��0����OK����H1h'J�Z����E|�(_A|��~���'"�*P�D@;�YP�9�q�a8Ȏ<�ǧ�G~Y�6���nlfy2c�5$M���"EQ@����SL$U�~����.���8|�"'K4S�e�^����} B��r�#�@@���727��TX @
� 5�e���H�Ͱ�n��L`'��&bm��*�䐼2�+�k�o�&�]$�jk�<Cܹ�>]S���Hi��ڤ)#�#��mhc^[Y�Yk�r6�T�dd���R��(�j�j�BE�ّ������@�<������3&�A�R6^n����qR<����.�����Z�/ow,*@����*�7.	n���v&�P��c$�(.ݴ�)����'�>�<X!�W��N�j22��\(k%K�V��'1�EP�����[7�Ɉ�z!yG�dH�
#
!�rʅ�{	��GJ,�e�� �Yn�R)����(�bh�^̳fV�0��nR�MB��VP2lJ$_-NN�D��z��0 �1�ᰊ̊�� �3��៫pN��¹ s��l�: AMe ��y�o�3��A_/=H�����ꂉ �"2!J�
��N\@�X�M��/ȹ��D�ͻ���	�|�!�I�G��`���J�?`E��@��H3W"�NF$�
��?%l���
V0�Fҭ	ԪHE��
<Hc��Y�V,���".�b�x��(���<�P(K���l�%#�Zr(���Z�������t�`�c�� ��?�˷}S�$w7C� ��6G05� q��ƍ�����Ar��0a'��/ma	C��N��͊L�J�d��G? U��K�"m��Kj�.R�U30���ng-̌�{�w��RpC�^D�ot�P�=ؙ������ C��'��?I�wJH����z��Rr�h׽��!��#�R�h��B��{!�]&^e,������07���C��,T|k�����e�Õ�5~N��D�"m9Iw�:c� �����Q�@��*H ��bf�\�ce���'��T	�5E�����ߟ���j���������۫*�ł�76��T�UAnn�"�~j.k�}�r4|lG�u����tT|q�ݎ�4i�7_�1�\Y�O`$�UӦ�Z9X�2����k��f��r�G;J�B��f�$⎣]
�ɡ3r���\(0!I#'[!B�+�L�����u&P0�T�E��.�!L��?��Ȁ2Acb�E�����*P�{rmոH*Q�37$3�� *k���\0\&�j�6��\��v��Ԡb�,аQ\AK	`Dc��Q����441#����ğ�i���I��r�f�UWtg � O�vD"Z688 6?�KQ���jF�<Q�:�FsZt�������\���Y���J^\�זD@���B8��a��!�{~�܃9��rv�ølxE�5�9�R6��A^�uk�a�Zǣ{^�_�t�����r��2+��ƣ�/Sg����3���P��:klf/*�z4�o�\�YE��˘б�ݫt@u1��!`q ��~�2{@�\�IKv	��h�H��YA�{�`�Z\���e�<p��k'Ti��h�`�d
�#&�g����fy��?D�9��Fi��5�j6�9g,ښ������ql6�BNX�'D���Z�BC�[|�6btń	XDY��Ɠ��J#����눹=��d�c��yz;�+^��)�E��&H8�J��O��ț;m=�B���lf�P�%�ȣó�n>}^Ҵ�qZ�D�P�Νj+k���4{��x���-hF΅dK
�E�2���X��kѧ**[:�PbN2�����s������6~%�C�x�S��7�����8�?B>��4"2�"���~��	�ڑ+}�\.A�Y�LG�5S�zT�sE�N�\���% B&EG�Q������u"?z�����0�㻠��sI~Jo�9;���ʈ˫U㪌���o&�q��2�	�{�^���(��_�ꨭa�Pc'������Z_g�i59Y�Uv�����C�c&n�#�l���*%>����?+�7��{_����N�/��z�s�#p��k�y{��tob��917A����|�#���ٯ{��Gz=���tTtv�����7����߶����Rw���͈�������?zh���ڜ�X�k�{�����N��55Z4\B�����Ѵ>)�o��sj'�g��s��ھf��W�'�Wd��F6G]�� +���_)�k+�N�2�U��L8Z�r�"(���\�ƵK�I�vI �7���x|�LT$�Ѳ+���@�G�����Q����k��2��?'W�~|�؍m���j]El��7��FP�5k���*�/+^Ȧ�gz�7�- ��(ڵ\�D��g8D(�"?ro�U ���~�D_������q������{i��4ظ�_*?7�6f�.��Ԇf�ⶽ�Hf��w�Vx��� �F��26t�/9kl���m؇�Ƥ=�bD,���Bd}���_|��K|x�Ƀi�x��??�|c4b����t�/���ߤ�E��%���$�'�\uJX���&�&�id7� D!����xQg"��[X�Q����S[[KN������\F؜sX�>m��`�n��(��vAcJѺf�0o�r��2H�uΑ�\�6�����˥f�9c��i��V�H��)uEk��L�ؠNO�kLF��7+�a�W�� ]�����Yƺ�F��nI���{��H��}�w���������G7CDA=��>��`�5 �ܣ�m-�x�5�c�c|_IgH;,�洌�� ����0x|T�&�/�9oq7����|n?Z�fz�l\�%�|+5TE{���_G����#M$�Oh)q��w�$�]M����g�쏽S_\�TY�4�#-U�ݠ�6}�r`���`��s tc��2�%����5�����]�ק��4��L�mz�!�����"V}�N��d�2���1G\���ޙA�o�@�9 �i��3��Y�NYXQ2�-r�m�\�i'G5�|�p�d��Й|�GM��I>m�I�"Х.�kD"�m�P=ƁV�W*�v�|3���~���}I��cp21Y,b���!�ˊ@Â�h�o�.'ZM�u��17:RE��XͥQ�j1��<����4�?_�<������o���3�ϸ�  �8��߂0�|�*Rc< _R~EH�j�D��׹\<�k�UZ��U�F>��``e�I�Y}.��/�������ퟴD@�*�*�t�_w��G=��:���NgRkd�q��qyUz�gh��M��a�#ZC��_���W���鎵����ɻ�5$��|�m|�A1*����&+!ҺU?9���]��7� �������x]�A(�6�$�V�1����5�O[�h]�F�`"*�a �	b"1
 2k���^�t���U�|, s.�j��Z�Ty������LI��L�>�s*s���O	��S�?��}Q�����n��z.����L�b�9&��� ���}�|��yN |��=��{/��0�~G��-z�'���޿�s*�����@�~���<y��h�}Ϥﹾ;��DC���� �����������T���˯���d" �A�� �8
!��EMj�7#�!a
�1B�A]5�T�4����e���"$/�h����@!&�(��FO����Ar�a�D��ĕBH�R�Cbc����[��d��L�Ex�zDDE�.#Ɍ*��A�d��	�|�%'���|�N@�R��ZD1�(e�� J�0x z@�_��E����-�}���P����d��ɟE��>�����,��:|�|g͛ b|T�~�M���M�8�%}�K�>}+��k>a�Y�Bu��l
e�R{3s��1�3dF�ɪ���b?K>@)>����n{7	�HMY�-D� e�d9�����C��>�!�lˆZϨ��W~X6ga�b0Y=4�,-mْ�j�.0:ݩ���� 3�$4M��i��|������,F�Bb`ƫ��U� ��4���/�ftybnd���'(�wH��>����0�-N��wF0�H	�����݌�7M�Cf��S
����R6#`�),�.ݒ�ki�G��=n��f̀Ŭvi���V&߷&L�$Ϲ2BHI�92f~��/��A~eW�$�X�[�}���2x��\$�Y�'�+��N�u��6E��HI9�JH��@&�H�+ۻ�"J�A�|�~I�n�RC��RȺ��!t*S)�����*FE�����%Zw��z߯_��W��)Ż%7|M:B���E��̘3���edT+F��H�IDXMB9R�wN��]ɋ
P�G&ɻ�.%4�u�1�$�NN\�8j�-T!���&¦`���PA,-�.�j͍3��b��(f�� ŉ��{�u#׸�c�><e87o��0[��J
!�u;Z�Uˇ' d!#V[�B��.s.&��A��n�ɰ�A�	r��،QTL�U�SR(�*��q!\�4L���$[ �8��]���nژXj.q܅A�ۚ�F��̶SV��.J93�%3T��I�D�[,G�� �R�܉�x#Z����*��O`m���X��pY��[l�scɘ�1�-�sTNZ*��n�)�{�jS-�"D=ҜCH$�I�dY�^O+o|�Ԣ�6�8�.��s"d�37S&�2�%�Rm�he
�tER ����Ffґ�n��\FR�0⡻
��
 �J (�rB3�ȉ�f<Q�H̑*Xbg*̆�!�9�U��M�\�< y�O��"��@��ӊ�ET��LmZJ��[���Z�\���R- ͉6���"���b�Ջb����ВV$�co���o<����ңRm#j+��ŊJ�M�J#Y6�L6�[�h�dђ��3�PʌDd�5�7(�F�֙ci1>���]5�I�Y��p!���S H� "�W^˸�+�"�~���կ���-���e���!������GT(#���[��U��:��{�@
���@ �� �@0*�#�J���"�
 �0*@�B0��@����7�M���W=��o���w6q�7�Ɖ!�(�ġ����rW#���5�e�����;��E,�R��.?�n����'�����A��Q��?ogA���Z��d��"�j"2��2� + �H��*�� �	 H���q8�\^T�3�uͱޅT�Ma�*�歽��G��9q�v�.or<M��i�$%� �J�s����?��2�1�a`�	b@c9�|p-�-춸;\2@*��r*z����gs�랷�u�-�wO�������Y����|�+���s����}M�p��_LG����M�W���zؾ|���*>���|���\(�(����/�4���g�G֣��5�����}���O�䟚���ЕS�?�w��}��y\��c���;���L����y4���߿���O�_��8�������﯏�W��-�}����qy�����zOK���������Û����������#����H��c�<�}�|��Y��������/#�6������>����ٻ�c���)Ǽ����=���e��B�n�j��n�ߋ���?�|��6��ٻ��9/�{w:F،����|y{�g_����8y���W������_���y�U�ރ��^�͛�"�/<K]c���I���#N���Y�Q�ը��/`9b��x����������:.��]c�u�c��˳�^[���c���G��+!*�5���d������`�*���Qub+�t]'I��΋�x_2ϫ̟��)�a7?EV�k��/N����6lO���W�����/��~���U'�����zOI�|�&���t��[�կ,�/��n�Q�~p_�ܿ�nK��.�=_��x�.��^�?�+С�<�z��d�ޫ���K�����*z�	x�pM�<�͔�f	?��>Ε|߸6O!�h���&���I�����V�T�������~^�������h�{�}�����}����_�n�������<�����~^P�����yo@o�x�����%��^��m�}�O�t�KK�A�G�����s�����|���8<u^۾n�Mo*Fz�y]�c��sܶ��w�5��o=��6����G�j��=��o��,U�aG���`E	A@" T�E7N�������.���ь~P`��ߘL 	e�p��^E��G]�'�2���c�9����^yŌ"�u��Yd������W�Ȝ��C��m�P���v<��r� $C̱:��M���03-U�t�$�3�la��#�����e��������K�lfyi1�w�q��P0?��<Z��c8 1�� g�Qt˗剒X�XK���C���ɖ�y�!�b�X��>�vM��@�낟��x၁����K8�� `���Ս�_x�0䷔Ͽ#�U��S�_���|�Ҷ5__�& ��@c ,���plbCZ�X�t����i_����g�ܘ����dF%�x�\n �v���-��܎s�k�E�3���\C.�܃�0�@$Jrߤw����C�|6�Oa�Ǭy��o�_<�ѻd�;��S�F����M}|)���W(��E�ӏZ�=x�_Jz�ٚC�%Ͽ�r�+s�<��uM3�͙��`c�0�����\���s�3�q���s������w�����{ac���έ����wd ���0� `m%��Au���O��ui-�G?�I{O�4�ܗ�e��q��f��M�����3�c c<�H)1�Gc[�����n��� W��w��������؏�_VW��%����Q�p�~T/w��c ����k1v��\���$��b��,���|}�C���r��|e����nw��~������*aXt��O��X����׋7�˴��n�uhi��WBRF�����1�'/��$ 1���Ϣ�lY�W7(;�H�?}���K��c-�Xb����c�k_���v?zWϗ�~n���%���I�id���ɳ��ϫ���<�O��� ��0?d��c�ո�y��Hw���֬�9�c�}&����;�l�ߚFt�Ԡw7� 2��m��+�%y��<�����4��s~MV��������/.�!Ȼ�`��S˗˯.w�1����Q�U]e��Z�`Ϸ���#:���Q����h`� ɩ����Tn���3��j�����|�wOZ�5c�����}����i��g��0B߳��ϖ~C �`c���Ƚ�k���_=�p��̭���>����駁�)>=�(Z���<7We�?4��	V,/���۰c y���t�r��m�ށ��^Z˖���1z�%��� �fG?/��`�f��)����x F�xm�� 
ߡ|�{���;����,`cr�!������-IB���ӟ�ڻ��vn��)�����a��u�)Dzﳰ��H.�^%�)�j��}�����6����ڕrs���9�����FT��Y��S`�1���g�["�kd�Cgz���1����\v����#�/�# `c��S�G#����(��ke����so�Ε��_�����]��������ɝ�=�vm���խ����>N��>�����{z��2�2� �u=Ϩ``ct��Z�g�tȋ��=|��CN�C��ps oʿH1�c�6���c��ܼ��R���}O�4l}��/KE�k���������%��~_j���g���g��W��xO��j��D�<�cP�]������u������ӷO� 0{_�ƘO����7�Y�҈�d;~��w��/>s���p��Y1��uz��=�L�~�y�����o}��F3��6�{���+}NX�U)Ϫi���|���7mW����J�'�䴻����8}�˘�QKK���~~9BXI@01���B~:�\��W�r�%ڏ�V��3��c����Zk���|�n.� c�W�>��%)���QL���G�T���?e;Xo�ٌd3>�yu�ь M�,�f�����`����h���
�Iwٯ���;���X�:��fBQ�*��߲	ef0_*�r%η}���KD�)��N�Y����4��,`���c `��������E�r˧�wHӧj�)؅�~��8���/��^�x��#�ٴ`c>y��j���v�}��:�k��o�\�,���I��KR��w �c ��eaf�-[�=.�|�@�m����ߦ�x��~�FYJ�B���/�q���xc!��?��C(2�~�O,kĴ����k͌�t��?F���8��:1�`��ѡ���#��WDǦ"�z����Sʨ�01�cϐ��Ϫ;#�i�����l��!�}�]��{������|�>_]����[W2�*�M��`���``d"2O�޾:��k�q_Rؽ"����w���}z������>�	=���� `�o��b����m̧%@\�5�>���J�{�>�N),�ϒ����б������ �ܜ��Y�� �3���ŀ/�����MG)���Ew5�i�wٞ{�9�An������w�Hy�w���9}��X���_�~�;BR���^�}��qC9�����R��3�y�zz*��Tq-\��=m��'�$���=�� 2D����BȂ�[�]��;]���~~�>�D����͹n���0�����m�;�uܷ/3z���ف�ó�ĵ��5�sY@2=��!��#�h `�y�����T휗y��I"�MC�tP�휦��俁f��/���c `���6U�p��Ռ��ꏽ��W�TT������A�J?<1����M[�tE��%���c�����֮���z{O[{�[N�O�F1��"�Yæ�_����/b����N��ۛ c�>�	�����5��Y�xX�i�}��n�Q~���o���tT˾�c���o�5��bP���0���ZC�>�v���M�C�~N�<M޼Yc�����|�1�1�``[&8Yu� ��8¼�������eF1�8�Q�Z��&��j�X2M��'J `y�Ov[Ј	t����c�'�N徲��ؐ%R̤�
f& �fؗYIg4�H��Y=���Bl$8t�d�Y�0�6G$s��3�L���"N��"l �!7��F�$� �a��E+��RVR�!.�!�c�0�ZB��H��^=��}$�͚c<�5�Z����� �L��+��M8y��%H�
"��:�OWO\��ɒVw��0�vr�'�IXd/)<`zzq`�e�\��FS)�v\�$�iq%�rۺGkv�X��,\�����h�V20S������.��B�(���
���8Hwn�\!��l�����,:��ٰ�r"H����� �ݓd
l��'	�02,0�D0�;��B#"iIGm�C��s���,�i2�֝�]�Q ��`F�ݤԂ���e�q�#
ڬ-�{7���x��i�$c��F1�m$�`Q�ʈԆU, �f�p���m��ʑX�Ee���u%�'3�!c���;)�ŗl&�wN��!��$5��m�#K�5�,��7J�p�JS�JH�5�p�0�GL�f�:%͚XK�l�iK��B�.���4ʨV
�\yL����io_�bD��ՌX� �+wA��d��e�N!v鉼ێo=����X�oFq�� �qY���e��r�@��(T�5��J�k�;�'rB��]��@�m�$.�uYvЁ�1iU4{��H�0�kL��^�.�1��a1ҔO�Ri4�:b͗N;�Yxa�vR���
�TL��V����ۍ1F�x�'�l��R&�H�D�WG��*5k[2��5H��T�1"s����;IZJNF'(k�Ԋ�h�ݹe�@ĉ��"Zf�DK�
f�c0	Ja�T�R�[|��9HC8	�su`�����]XC4��o�� AdҤ��K��g1��c(�Xk���i-7�5�:0!a�6�(�͌�YĦ��8f��N(az�:���@��"ąd���3m�&a���ouqa�k4�����w\�r�m�	� �rv����1ik���w��d��n���h�-y��@�&F���v)� �l�]�d�	�D��'*��0�R��P��wׂ]�w`	@�YL&�l2�!e�l�$&�u�_l�퇶�rH	���ݴΔ�ꐖ���DAe(s"slBs�l�8w.씄7���vx� J�$t�9�,Ie��<o:���u�f�z�r��n���=��0}��7Ik)4°�f�� ��1�4�g^ ���YU���{	I���n'^�]����a�UۚXGalV$F�ZK�9�Lޱ��z�S	�U)-;i4�Q�H�zH���t��HA)�ޕa"o2ul"̏c����)�v�E[	������]��0EBk��=f��픐��01JJJB�+Vi7���!YJ���ܲ�d4�3۲�����۪Ȝ�,ݳ(�n�z����:���)N^���k����H�#���Mmv��V��VD���b�rl�)m���i	ZK(��2���ll��
Ջ{e,A�m�N\��ٺX��I�5�E�8oZB2W���e�� F\dL�J^I��%�i)t`� ���QPu�]�R�B��p���p׍ C��� ���Ȭ��O2�),2�BL�\7=R�Z	 `j��i�|f�o��Fq�0�Y���B�To=ӕ�`}$�[��=�gi�Ô:q��z��L�.�u�W�d��S5�a�g4�̓=�B	���,��EQ7`���*:|o�m�ٗ�c�Q"��	�&+�PiE�B�T�34�V��i-A��%�[#9L�P��L$�dA�u��gn���T��^X M�x���q��Wͩ��2��4	���l4h�)��ѻi0�*<JT�,�+2�UL�-1�5��e-b��j�wh�q���SQ%ݞ5�����sM
2x���kHa)Y��ňp
RڋTli.V����`[i�uf��٠1_e�v!V�k7M��Ê,�`i�lH-TH���Y��_ � ���`�̪��2����Y�l��R�fL���3�H�	čQ�=�vs����D2<���e���z�m����H]���Kcij�Xw���l�B�
om� ��ӝ��ʯzX��C�$��KM��5����	d`$*B�x��4����T�ZYpB[+̳^���t\0� h�� Mځ�4�3F��M=�v"g�H��Ą��6�6*;RP0(έ��)4�k}���pҘ�c�gk���Ik-�T�`�l$�Ie"C�i)��ya�c8�,ư��k�鑖{�xKYy�5}�8�("$)KD�aMJǘ��ړJi.�5�pn�u	�b�yilbR��M�+#F8D����	bm���gKՃ�����)�/�f8@�#��%_� �R�m���s[\`��bė���a=:��u���:�m9�Zu���F�o�i�V@dA���`:�Of�l�����OfG�f�@BU�fI&�0�
�̰�!Tiii����S3)J��A0*H"0��Z�Z���J�V��!�,���J�z����,���aa-�I����'t�4�a���)5|���{K���H�l��4��C]x�����c� k��YOA��2n����w�]��O:�	�C��ZBk*R�a�)la g�H1�-Jx��qP�����|[�kj,��!�l����4��jŌ`�7�e�1�C]�vǶؚc@P��#4�A&�Q^c �4j��*y�Ju�gN�Bx���#�Q��0$�e!J@2n��ytb�t����zy�׽��F�̠d}޻�m�N�*ᄭ��!��L�.�wj4%k�.Xi$+���K՜bk�bN�|�XG\���KUaR%�o�Ҏ���p2Ō^��ե&�����;��3I���M�w��:k�R>+�/r@��0��__o�>CU%�V�F�4�@dB,2 �<4�Yj�op�m�ܲ����!�'8BR&i"���p�x��-�[�v�l�6�1����#�<�'Q%��@�-�K鶓L��0'o(�>2��
��ޭu��wY�aaz�$EU�Cn�ṪX���T��)��ĥF#Pu�g�Q)�&�����`:�@ �$�:	�H0Zzu��hC ������%��kݳ^�3��Kl��"aI嗖�1E0�&�0��2� U�s�Z�iI�3�(mɰ��JP��@�ik���	n*��|f�p���XH )��a9�t���&�T4��٢RÔaP,�� �b �,���a"��ݖV@�WFU/v�r�%���%�0V�Z��Yb�Yc�w��Wvz��7SF JR�X\YS�&���	�7�應a%"a�:��>S(AU��_2R^bbdB�n	��a��H�8�۠*�|K�W�����{{Y:���w޽#��T�xf�&i��j6>�7gRη	OY�^B! u-�%��f���j U��떹[b6�L��­:41M�v�v��wo�f���s;��)$��)h���D��*rԊE��{}�ɦFSZء�� Ij! ��Cn\�G6�m�10¨��mVi,�&[utr�}=��� xJ�(�h�,���V$S#
���cn�,&��4@β�F���Z`7 �	��n ��c�.i���\Q ��$G�b�b.����3���3�)��Y4"1�\Q�G}�\�q��Z��,���=�[׉u*��b^퉲B�4���q�b�9Lb��8IFU`��(� ���$=��;�0"1XC���(F#V[0pA���5���Me��0��B7�4�H�K�� 4���v۾x�&�V>Y�@�צ�RR#�7c@B,N�ml�i���l�0��0�^� Ƞ�+Y��u��,ke��l�$��:�펱��UG��1������ݎ�u�N�K�޻��R�m�3����#XBѵ� �^=��gO]�+XW��͕��! ��c�#Y)�펁!��PbB H����OCI�GYHe�회�Z��uF6�%��G��I��l���@T��s�"2�4���2�!q������ou��n��s��q�B�f���&�h�����t݌��P#�7�nФ�f�L�@�8@I�mL		}�]0��0�yd픀Z���D��Ƥ'u�a	�D�S
I�Y̖�m	Dy�Y��e@i,�N�����l�
@l�γv�m6R�S]݀M�I��Մ8C�[Iѵ�EU�m����k�MdڛF�X���r�kI7vhj�<i��q�\	$k�jCHz����3�nބ��"+"$L^�Dˮ&n�\��"a/X�6�m`,�4��ђ�	����L�X#�\�Èɰ���3��6�rx���Kd�<�,�2�P�i5�X�0��'6r�5z[7X�,&�a�1X�-T��[����С�I�Uƨi�r4��'s��'W@$�2SjJ�Z�:�EHKb��֔�I
�P'�=�I�<[�xģ�W�dr�]0�R1X�5�ցdI+&�e C�U�ŀ*�a�7c�cPV���9;XQa�dI:�`E��2�wl�l M������lk���T��
��h��nzM�
A��뤔ՌT��i:���^rK��X*� F	&�sd2�)ݼ@Ԃ�@���k�$jW@��@2��B $Ci��!n�Y� ƋeH]��Mv�"Z�N���o;X�
F,�4$%��e%�e�;n�BQۅf�,Bb2��>�Т!��-�ZL����&�U�v�CX�=E�u�k�n�3�ɰ&�c%��v�wM�E�Y��6P	<�⊬���+���)I@�,�QBP��1��)���Y\B::�&�K� !�yK1׷IVi����q{eΆM!�\��O�(���6�V�B���lk�+��,�9b�S'��#Q����RQPŚ�M��D���%�mn���B���S�<�D����uaH�X�"�q!
$W�a�;x��.�%�F+�yjDw2%!6=R��Ƕ�!��),�bD�fP�*p'R�A�XR@��Nf�Y� �L R�^#U$�U�rk)��v�� �m�t�i�lg=`Պ ��P��C��6��b)5B{��E�O�E!�OZl�L��3��!e����u�l��ݩ$
uy"�M7�ň�!XF�gs�z�\S0��_7<�b�)H�/[�렸Ddee���V�b��a)-�)�q�i��Z�l&���`@�k.�mo�
v�Zf봕%���g�D�"�IJ)�P!J
v�
 "bTP�d�� DOz!`Rj�� ��'�~���g����e�߹�9���k웞��x��������w���ɲ�,���s�j�����m�u�����/�*'X��J� ~\��������akԶ1#�Sêt���C��'��#�*��)��Av�g�+�&~�Cq���a����4tM�H�sa$2̀ s���q"��� �p;��� 5���k`��m�6�F-`3s(�����k�U8^��A����f��u>9��k�!�fV����F!vK9�7��o�:��+�(����ErUQǝ
��H���Iw.�[ߘL�N(o|e�RI�^�J���!֡u�f����9�&px@��J���8(d�*A�H� ĳ�@QDЖ�����y.��s7���ڄ�d<�l>Q%���V�U=ZU�5�݂�'L��!S����Yb�E�X�N�j�RJ��\r��v`^u$�[*�b��w�B5p;S�i����TX4x�Ay�Yu��&i��n�!ˋ
:�>�!��ҽS���P�[�$|�G��x8][$$�U��T�wm����(�&5�e@U�,��q�5e&X%��\�=|�̑q�d�ƌz��gwE2)sӆ'L��πY .�
!�X�r��*���ҳ�n�"�Ge^��������Few�,�����"�P�;���D�	5�!V��B"1�����j�lr����-WgV]��L��X��\�i� s���BI��A��� �\q�`��i���,�FD��Gf�����l�%��O�a���C�@^a���ϑd��V
���	�b�m�ם�����C�H��˴3j��n5�jr�qN�t$?�" ��د;Vr�]�:\�(ǹ��V�0Cgq�W!�C.m������K�[�Y\��oD��y�K�'�P��x)=ċ�x��L?���DK�l�Kͯm�qk�Ԇ�ͨ=���,���T�4f��9�jY�&��`:z��"+Yp�^BAč�2:�3�gn�3߼���2�&���6����R���A�QLĶ�(M�f���iS'2��D%�̚��Hv^6o��n���7��-e$�d����&X���`Z��0��~�f�	�.J�A4�6��A��&���W�٥�%�WAE�C�G�����
��I}k�������[��X60�|�)Ƈ:vװ�+Rg"�u��P��ɀ/�g��[e�Y�f�����2��]��O+њ]�ҴS1��opl>>���in��@�T��s[�geAS���=仅�Z��/k�D���Z�~���V"�b��FY,�D_H)ĊX�D��(�"���E��CDJf�
�`Bd�_-�O��>���?k��_��?�Om��<���fp2���=x�z,�f[���UMb�aw�W<a�O�:/����I�I�|8���ץ�?]r�,e���[�����N���Bx��'�}��#�$��\�6�!��6r�c_�ڂ�����l'r���4,eA����@��x�~r�XD��7�y�2%9
x)O�!E�%��b6dn`m
�V����.���$�rK�E|�����,bz��,mF �S�-�r&L1D�؂�fXy�kٶs�\Ԗ��ӓ42�(S�-�f���$㝻����J-�݉�*\x�@x�61l�8���@�EaD�;a��@��/��0QSltJc��f��sF��&,�y�*c���D��(�pQ.������Zk�ҧ���bY����Q�&�&��;���T�I҃�*8T��F�g�=JY����u';�ǋ�2�i�3Di�i ��fJ�bFZt��ϜrK�Gg�)��=<����"W�V�<
�;;K%�S E6�Rh�,P��S6���n|����`��\kzɵ��}�q����83�<��(.撁�
��]n&�Q�5i�¨`#���Z�7��c��RPRKL���wh�v�B�̹M���ӆh�䰒��.X�𭋘FdoZ�n%t�Yzz�d��х!��X������AV���!w���TlI&�j��b��$�eT%ܮ5V�z�mI���b���lN���T�w>D�
[ҳœ+,\j�R��-ZQa�V����!)���
<�m�O����z����$��C"$�7�ޫ�`����<Ӫ�V�8�P���M�e=��g���2�"��R7���8�H@?��Z��L�iH�1Y�FO�B�}����ݚ"����<�2B�[��.Ђ �h�氢�7v�x�Vs�b?A��+lj�-MMUrCz�[+�q*w�8���i7�4�;��@-M�L���ې��I-�x��!E�QR���P�۟`��2�6�ф�DR;��l�C��W��	gl<O�A-ͥ1�����b�
ar�+(�������pL�z�P�$�0p���Qr��lt;!X!$�	0��� �F��ͼ��޻��\�)s. �d������u��hp+��������	f4,M֥R��!����(�&�̳��CO�:�ީ�V�`�H o�2D��.W:����!��������[n	H8�� �([���i�L�a��-����b�zt:"�f����t@=Z�� �U�$�t��0$��`k���a
Oyd�Km<��ں�|G暩"
��� �y����ui�#�3)���!�p��Y�\�kM�l�5I�EI����o#�6h��)YU��M�V�<�!u�e�����v>�h5)����[#���:�#��M�{dC�[Pk���O� :ʱ�#
�*�$Mp̚=nLS�A/b�䀶�?�C�c����RTٝ,1U'LL��t�nC�]�jI�Y��b]�jm�D�A�YZ�a�7��ht����)S�Gf�ͪH5��0�����A�Ŕ5��	&8ӑ����;o.g���(��J�$# *�"�2)�A�����%~�O��n��h�
�$`[#a0!�a��L���!s�K%r�y�e�c���0$\��by�<��:"�wn��BU��qEqJ$�L���:��p
�"!7Ў�=�4Y
*#	Q�1k!AM6ƀ؈э!�R2I�I&(��F���2��@it�������Kh��f���6&���X�1Z(
(�&��Qh�A[ѱ��&5�c4� �C� � �����F��m�&Ō�Hd�DVR�2�h�(�$I���&J-�[ɔ�(���Z0j���A��	�))�I�h�F^y��-F֭"��8!H�X��!�0��}^ 2���+F�5kF���J�[��V�����ߥ��X��E�(�A�1�,m�1E4C2l�$Qh�M�0ZN�P��^�Ţ�m�Z���ڹ]��6)��bƍcZ��\�s[�(�+�F�6�.j����R^Z�^�54�HK*D�@IK��bE@�)
NN�Bs�ϠvA:��;�F�p]Bd��FB�$R ˞G�2�
呩]hf����4M�qR��%*�I(PܖzS&�i�,��[m_�uթ�w]�mn�<���C���9NG ��4�sZ���u`�C�5`L�X��Q��L�dBe(f9���!�)��N*�d����PP4A�� &8����f�u�\�SM�
�At����+�����BN>nY!�E�J+J�"��E��j�Q|uw��3i�h��mk�D�j�P!4�J(�
"d�i�6��鵹o��H&@�y
Jr���`$��TN�8h�@:d!M�x���2��� sL`!�(2�Id�PK�&I�6�7v�p��#��$�"���	�(h�o�AM�*���<C L��hh 6#س@� ;�+Ǡ/	: C�~XW��<p2���*���H� �"����u�<!G�Mǆ���C��A4.0�Cl9\���� ���/y�h.��f!�&bG��(9	pUN숩��y8\$��Ƙ0��	�9b&C!G��h�J��u�h��ѣ�ř�&�{��լjF��&H��p�� ������'�Ϯxo]�'�>O`��`����]���6~�=���`̀���������aw�ܟ��W�y��mr�0`��8�4�}\�ߧ��
��
Zy^'��99����i�I#���|��������f�.�x9@!��O��	f�)S0�J��:�*J�h���/^WB �4+����|G��
��&uc��FJ!IB��O�l��u4 )0���$�����V5e����h�Bg�r���:���ρ�����qCv%)]�Q�������S����)�W��������I��AT�)&���u1�m��Աoª�`"G9�AJ��YJ`%^J��RTԲY6�j�d9F|� s!��`a�  bSb��ݲ��Y,ȍ�Ej�-�On�QIoun��%J`�1,@D�:��!��H
�R&pj�$� ��֫\��J�] ڵ�2�-I%����ݨ��ۘ�����l�K��k��3&�k�ɲ����̳��v^5v��ն��5�	S#$D��rD"EW@0P��G�@�(�!$D��	 ����%AU%QDH �ą"�B6���I���uu�d��UU+K&�R�D�F
��H ���B��* D̵0�IH�9��U=�&B
ʫ@-�H"�(R����i���z��H�?��y��^A���P�fL� C��ι+n8��û"N��YX,N$ҁ��9��D�뙌4�-�͹l�d:FQ���P��T
;E�h�k���Z��H��B��Bg'�jג�睂�5Uu�(�l�3��́�X\��)�a�ks3JL�J)� ��QS��"��T�H��D�ś��i������tٹ�&r�6o�,�|���iEaF�?F��Л(����`۴T�7呚k���K����]�3㻥��/��;��S��HݚCf��ݝ�oz�&��`r��]��,k��WϨg\I�+y�eN��r�v�Ķ[J�ޯ;�'�͎#�p�������1�R��T�)u�\<iD�ld��q��u��.Ok|��HRvq��m��˻ݗ�N�<N���x�PI�XP�� ���ެ�ݶo��3��9�u�z2X��֤-&�ݴ�5���Fk�[�i 5VoYhH,:�c-��d���i�m����!��3�i�[7A:˳�l*��۴3}��vN���s�+5��k;��6�ce��gwvlH��LJK�	R ��i=�i���i滷}�Ug���M!����66S(�)��	<�QyJi�]2��a"O	Mc4�<u���ư.M_o��{;w��rMH�۔ʲs�K��q���8�$��$��4�EH�K̳u�<����Q���zy�������B^��9��KE���}��{�fԈ� u�BV>24��B"N|wN �6���!Ќbf���9��åc,�ia�`�!��,T�����λ&�qB*��D	5���j�ޯ=7 g]ӣ�4#�n��aN���4؈�)_-ݗ|�%"@}Rꚮ��4��N����h@�m�z�v�_j`E�Id=����Ne��2l4�o�hA�2�K;Z���aa4�nu��p��0yp�4�x���*��֨���D�͐]�Z�x�1{ږr���m�onl�lp����fXSY���\��%8�gM�vy�t#y�ӛ<� J���q"#���D�B�R8F6���	�sJ]%<�/��.���v�-�,���{��x�I��ti^�M�0G��V�ݲ���{���=ݽ,��Rv�!�KݷJ�i7�`��gK���i��c!a/8�@������ύ޹y�y���6��:��:����@�U�6������0#���N8���8;{Ea���ꔉ"�^L��'�V�&�Ki
���1<[[IM��	�/y�/]ݱ:��g����c=g�j�����������k��Đ��"C
�Sg���4�����q�6��L��! ��4�)��c��5h�X�9��%�4wg��;���$�撃۾�8��"d�=t/2���\u��t���X�٭��"b�G��7&�I4��V�v���	/�y�{���p !��{��5��	g3l�ڢ�a�v�4#�J�OYL��I�owy�ЄX�&B�z붤L��OR �C�M��R�6�l���k�,6F1����H�C*��/3u���$u����M4�e9�O4��}Wv_AX�@��6]K�m[0�%�V:����&ឬ��p҄��c40��iaJF�*FGݽ6k�ٺ�n��P(V[%�n�a,>vo�e�Sg	�	;��fݰbx�pca�녡a��z�f���CF���m=�J��댮��q��k���YJm�QT���#nٰ^���E����B�#d�v��� �cf��K���	|n�7b\B.e=c!	�I/8�-gX�z���t'��c!��
��p�K�����毝0����ݰe�M\'kVx�]2Z��[)����w���=��K�k=v�ŰiI'B�������O=�˼bK��CH�2z��Q'��#6���x�60
D���n�d[۵Ψ�[z��MQ�T��͆�#<�@�4�*�i�,d$u�¨H����+Z����Ą�`U	6�&R�n�B+ ��XJbc5�����-���ݳ@�Ye@�!��TnM�04���=y�)GT!@� �*�����m�^=wnm\�66���b��S-�=� �tɑ&L�H4Ȑ�sI������
�%� ���5� �2�S�������r�*
��bC\�bW\��r�IB9�y�m�r�V�m��ɵr����MR��8L�V��g#������+�Q��!�m1�ye��"-4���`�Zm}щ�TC�r��k|�9` ��(� ���ȱ%� �/�0�EDd�M066LHF�6&Y2%�FM䣐�z9�:�vL}BN���ì��W��,���#<�t�L�����5�-}[��j��1�����=�������wt�������,7��\9rJ^qD�i���>���u{_������:�����9�� z����G�oy�ڀ������	�|�+��w���C��:�O��s��������}�?�=�����}�����?F�9�X��@�z8S��/���z��`�=���9<�'���	��M;�����| �	�9�N�B������=r.�eA���]�|�B=8�#��n��`���2�:����ե-V���$\���-����9ڎ�3��x�	b!5G��
�A	*P�G�q�-OZh�+�,j3����i�=�n'9�GǇ��ǟke~�o<�p���P����Ѷ��];�Uό��]U��҉?U�'ǣ���;7wap~ T��.0���I��3�`#�5�L�iD�}�mdĐ��'M�z�$.�4�g�0���'��&�%�(n��駖��Og�G�Ɇ���^z�Yc���&+�2�O�i�}L���~�K��D~w}���zu>�.��ܸ��vj�qdu�"�����t/�ߚAݯ�Mye�'-�5����|k��k֣���hN��\&���&���5���鵼;�k���+����c/��m��m��\�s�9׍MXS��z��kV8��}$�to�m���|��<Eu�.�nx�w�_�|d��8s�/�fx.���za�N{c�hi�鿿*/���N_�^����ˡ�3����2��\=|>�'�~]��3�/]��5���}){m�3�ˮ�ӎ�0�xCWAc�c>���-*��z�O��.�5)�a�O^�˹R�uwT�������{$��6`Ϊ
������3��\;X�����p2u`C��U9� )Q� B�QiU�@ *��Em��m����b�R�F�Q� D�"�"�� �����B��jՊ��c����bs��DH$���>��~�orC �]��s����E��� f���gNO���|���I� �6�4�H��*�Y��TD�d��+Y��X2(��Q��|�H]���IȻjM����km4���"�C\�WV2��;rjvF��t�Z2�QT�;2�kn\�r�@����遁1��I@�3dY�ߩ�O��d�3{.i #{K�d��vD9K2��Xcf����$Y	ݗ'ԛ��$�k�05a���^s>���!���5@�MG��y�%�W5ʋr��;�1g�>y��A�s�����/��XJPKӃ�B�2 L�"2�V9)���h�uۈ����y���P���(�� ���/
3�x���k�����ك�q��	o��������k�<�ogJ�}_9�FG��,�d�S�wu��X��ڜB�ɍ1��}� o�\���Pe	�5Ƽ�%��$�b+�)�u���\ݖd��u\�;�\�nE��^���[�Ls����|�Pl���{z���DƑ&[��U��<�\����O���S9i� �8)U�	Bk��9N��(1.i�	���9�<�v}�w��F]u��n���ۻ��LSί'�]1!�x�tԔ�0U�w��y���{��k�����[��l�'��|��S�<�?�@�UC������+��|���C�Gg��c%�d��^��~���b��N��s������.�����z�
�z�/TC
u�xS����K���/�w�nm%�wS/���4Cd�*\!�gk��>�ι�H�I)630����UY��M�#D  0�'�*�1.���#����|�/8��w�~��od�FD��RT�fU�����cb}T�ׅ�Ϳ)y�#}�o��t�}<��.,0��4��ݜ��nt݃���y~��׸��StX�C��2�K���6�rƪ�W���=^�s�ԉ���2i4���Fnv)�r��h%&�A��~��of���5����G+����R<�5�-�[k�מZ��m]���;�D1�柢VX`�Ņ��"��{�@Q�&�/u˻�1�˙&6��"� .~2�Z�{7��M�X .�A 0����w	(�v�$�S���-�*f�ǋ�+�;|a����[�jt��n���C�ֲ�M�������h�A�8w���i;�}H+�av1�Fa���z�o��K~z��.�@׋-w�Ď`�� 8���Z�C�y�	��Φ����<քk�w�y�ܦ�Ĺ�3T`���īm��p�Z%�4Hi�楧˫�ts"�]?�Dr��|2�E��}=M�,Y��9�������������"l&�±�u����:v�Y��E�˶�����/�ڔl��x7_J\),`Z�8ځֳ1ǁ��	.��XmV�w�+r�n���B8^A^e�}�WSYZ�!#����ֽd�.%��s~��4'���v�UJO��-�I�Vʏ�D�2�q��	Y�`㞈�t+g4�6���<�ہ�Z<�p{��:(�'y Ρ�S��-��H���4S d��	�.*o�<�$^�8�����7��*'����1�yY=B㖖$Jf�Q��^��uW�r��
����3���\d��-��ϔ�V_+0��a�t��I^x���,ؚ��L�ʢVj�9���B�+0�P:u���Q<��7��:����}K8���ݭ�R�,�-r�uB�����ͤ�G��:�3��L��df�+���|���!Xptfn%9��Z��67I⠣���1�KJ��Ñr[�36�a�Vk��^�g^��\�2�pW���D���L[���=�����s`>�Vݼ���RC�����@&2q�q{i��I��[��4����dj�wl�RE��a�#�Igb�U^/�=GlSM�7�Kyr�<F-}
'.��w*��t�B��0V���O:�jp�dI����!|:�7:&��@A=װ?6p�5�ˮc�%|�c����GO[R�G�K���v��d��x�3<`z�ԩ%�`�4��I�>�i4a�H���{�g[[ސ7�׺\n��(#@���+[�[��lOA �҅�p���F0Ac�'&x��V�8��u�z�"��F,G���@�i�6�o�(��VA>��po%�@�60��v�����]H`�i4�TU2����e��k�Z[C��A�������\�jJ�hU:l=���Qg-�f��A�,�-���4Nrga��,IV9b�J蹼,��ɑ(P��;�H+m,�"K�����J�\"0�pP�ɹ���|'�"�	kg�65��b�t�*M%�'�9vQ���Ҋ�����N\�o�A�3���*������Hj=���!ok��n�d�rH~\*�u�+I���8uu��kP��}�>cB�d7PSx���T�<Ji�3��k��.������a�&"#@�����Pf�]�ߧ5���W��*HSp�N�*�T�B#��/�����  x� -�`0� Aw /c}!�q	ܥ���-�N�	2Jf3����~nI�@��$��+��y:F&Ww/��/K�Dҗ����$�(�9���b���wX�W>Z��y��2Z�=�+��E�:@�#�E5e�*j�4ń)O�W|'��$��#>z��^<o3�+�f�����ҽ��Q�lx���(��BV-AG�]ݪ涋k�j��k�M뺸2�A)�p��㬏ezy���(��u�Ԙ��-��ȃoK���ʠZ%��(E�(��~�����6��)���g˥&��	I�Lhd�I4�HW-͉>����=z����g��k{�s_WJ�4J�&�@w4Ӄ��F*d��K�t#Ν�H�H��}<}oW&$�nh�F�5͌ccX�m|���-�U�F�����yt��wF�v_.B& �_���&di@�C۸�wk������� �P��:�i�����}i�h���ޑ��O���*
0�� ye�l3�x��o�߉��CQD_��O��/�2 �
(�Yc�$������f.B��\D#�'����zC�ߊ?�O�#��j���� xd/��MƐ=�@
��&햦,�H���C�& i��D�E��Af&��%T�O�e����%j�%��xE��HP I��)P:@rĈ�8Q��z
0č̢��kx���X�h@U�FF��H��Q ��ԅ8��ː�p��+%<0Ô&�	)����u�F�"�ńK�Y�x���>0��%�J�a�N+M�98����k�:�Dl6�xH(C�¡����@:ʤCՍ]�f��n[�r$ĝ��+C0�4��Sa��@�!�����\"�Ά�Y��euS�D�d�7fд��:��{;��@Ez��q�y����(ͥ�RFiD�Z(p���}al�2aG�،&����[�)���H.+ ���IB�����<��&��m4�v
�&�D1| ��ζ�O�9�#�P��:D���L�ڵ?t!�9�mL"\t�ɓ�$Pr{�&�p`�J#�� ���W���k��$_��Af�n�`[v�_.��� �D&r��f3ן8���p���P�m%j�"AMB5�I�;0��A�8�*W&� ��D��C Eh�@킐�$������=T�X�s�딗n�(�0������幨Y�'a-fr�e*��m�xA��K+{p�S-�:�"��ݦ��F�[-�'`�7� B^%D hq�댜$)���\K��M�TQH�tQ�N%�8"����,S�"4P�I����ËAq�����<lݦ��T�R+*B�!�9 7y�8f�rZ��Y+�H��,��QFN1DB�8�Z!DUҁ���ul8h[TbXM[5ݫXc��B����5�QR&	4��цB)�^�� V���!!o��:ܼ\�m���zLJr
�i!�@Ts�k�oS��1�'9a"��"�wp��s�ʢ���xJ2r; r�)��"�͹�d�R4G%���눑&"#h��OU�^+�*+�\ѣkץr�\� �\�Bn���}��NW��`Ȕ��[���,I�
6/����]y�%�a����\gu�竧wQ��\�3Ji0\��>� L�8~r4a�H�BL�@��b]���8S��x���Y��E��cX���o�mO���؁��M�@�4m�Y�Q�����h��O]�EDoK�Ƭ��_=���ou^+x�POwO]�1HS��'��\�j�&�t�X�����רBH���J㮌I�ܼ�F�7�sT
QE#B�%#�vi��y-���J���*�Y6��ޚ�-�[so�h�s���!��KQ�~�E�j���Kη6淥�[+��븃b�W�mnZ=�݅��Xۛ��u��n{e^"�(���׋E��u��q���u�E7u1-sqݻ$ܻ��i�8�]ݬ����M[�דj+���]-F�hG��$�2Kcrffb�fd&�x��j;���"�wwn�gw;�����Uwri���
��Y�+�`BbB �#�X20���&wS�wr�+���3���������Ӎ�m���:�1�(q�0c֘�����}������_�⻞��ٷ������/������<�;vA�~?��ar~�b�	��g�o��ZS����v�P�������
����'�ߟ�U?񪟳���셃���/����#��Mg6 ����H�RA?C��X��ƺ������@~M����F����5�[���P��{����;����u��?�o=?�a�gk�r��k>_Q�Ϸ�n��c���M<��{���}1�n�]����_[S�Pc������=��h6��s�y���o��i�g�IS�3��������#
~�,��~�?��/;�n)r#���&��/��z���(��Y���e����߷��g�g���]��������%�F�_vp��o/�v�k�c���]�����L��������.�������G1�g��W�i�7����	w wPK*��0�� =���.p��(F���E��k(Oz��F�A���^�0�g?�����w�$	������.�����?2�#A.tm�  l��W�}��W����D��j=s
}b�������@A�h7��5���l��&��%�5N1`������unZn��\+�t�+��f�m���E#��ș2I�C,U���]��MK��\�r���S��mz4
��ESEJ�%hW���{�DU���W�nm~Ix���|��h��ض*�{{.�4Hh����X��4[z��}���ǳ��Ӯ_\�6�W6�64mn묁�m�2X��o��^�߇mr6�Z��Z�l���B"�����c�7��l[^+oMi�׋I��rNW=wC� �4g��"=T!��+�q~\	�M�\H���U��vf�(����4��H�dܸO�}f�Z��^�m����x�� ��%�._ir�W"��Үj�cc{�C�"�K�	�Y�B��:@��Շ��Jv�>ϩ璄ƞ��Y������p���.����s��lk�j-Q���_j���Y M{-�E�ڍ�b�WЮVwm\��k��X�B�C9w-��zj��0Q4�K�5sW���7#Wҹ��J���)\�1-z���Q{+U�����,P��^1�wvy���#^8p#%H� g:�t����ˡ��bD�c��E�4ab,Y-:ޚ�5��lU�Z�ժ�|y�6�Fۙ�����^����sz�W!(M V�LH��@��9G\����	���\��PD*Wх�q��Rƍ@PE�*墴V6�]�9�r�RP�5 hQ³�ٽ��o@ǋ�l)q����QG�����깭��r��.�R�	������nb��9Ȩ|wL�D*#cI�r��|75BF(5����E�C\�2E�M1���f1Es�����D��t}^��h�$wz_Gz��R������^v��6�[ҷ���(m�;p g&���uK��Qrܾׯ^oJ�\M�5�R01Y�H�!
Da��'�(g!�	��0�$H��@�%r�ZQ۔݄�\���^��>6�h��ۚ���糡�F�H���^Jw�k����.��u�]����"��( w�T�P���m�|7�X׺ܹb�|-��:��\܏f��,�1�o���炙���&����oL��v�Y��F�V�����1 � 1*��n Rb!}>��V�M�Fܣh�Z>;��8���EI/gd�Ddј�MF�E��j���5�|�ً݁4���9ZW(>&	j�ș��d�8�8@���B}�����.��N���sE R���H����T�`TVv�xL������@�+�aWзyvܠ��o�]�+�>\�"@��d&0E3���b� ��]�sZ:��M!hhL�D��6��nR�so�7^71R���&.�(��+��;��]K�u�u�gnF��6��}�ڸ�� �r+���f�,�j�����j��Q���^���
��4[�wS��22gyy��w�$�7��	����]y�#-�r����Ug9H�%
��RȒ�m�h���܋x���X�xܢ���;s�#��M��$�9\�L���L�&]����nm}��U����Aޔ�(%�@Ġ�+����.Re%��4�Rk�+t�5��x��z��8��h�3/����^��wq�`�����c���B\~� B�~'߄�7�>�fXM�1Ue#�_e�� E�S�*	��	
Ҵ�(H����Z�R�h�6d"j4�-$Q�-	m&-�4F��IhJB��M+~����I������~�7���|L���i�O��5�}˖�z�>������|�"[�[�vߣش����F���gC����{&����_s���)����z?�_C��{�EఢՕ�{g���;Vx���+<E�Q��˷�QҨ:�)�Cwwd�#��. ܚGo��e@f�a���oU�����oҫ�|R���U/Nب��>���3��;�?�O�x~�O��i�VI�� ���؈�4����w� ��wp*�����J"�	�Sjר�Ѭ(�d�i-'��|y��+��H�K*��A�F�}���x��m���4�ԍ�O���zP�}�:��v�ST����`�t��$\���0a��e-�����	��$���Q�����t���l%8���ܸ�n\�B�W�8s����	F���ô���dd4��ox��e	SyZ���6���`I�(Gb�x�0ۋ��g3O��R�ePI&B�هr�~�󒖃��8�>��9����i�Y%Z;�D�J�_������w!I�qhh��*�،�����rUV�P%���q<�w�ri )���g��o5�4HzP�em��`�ԅ��&���%X���ը`�zv��/%s������<N�3׭��4Y�٢m�vD>��M�ݫj�䎹�{��L�����J�)N+F�w����>$+2���;����Vލ���4�m˭�'���:��|�O�K�wL�c��v�I���W������ÙN�����ˡ۷	 ��[i�ej��VS<��xHR%9��ϗ[9���ӎ@mK�A��~xp[�K�e���(8�+6����&��;06I��%4$���[2ݠ�/��/�iJ ��w@`�3�Az�kz`�"w���ү^X��)�/\�:������8�D\S/����c�s[�Q�6rL�U�ʓT
J�q}n�#Ӡ���r�&�]z��k5�8ui3�_u�ּܹ��4�(*���Qo&��V��I�h�V$s* �nN&*���-��35��
lwZ�|)v_&4�Dq�lg����N��X���x�Tw{��$����`�U�W�\6�yf��ۄ��w� b&����ʍר�%G˽]�,u�}�"����lr�g�����f�7m��X�{9�t�ǔ�:r]q��1g��5*(qS�60��A���[��4�gތ�7�@㣰\[�
��)]{?`Ң���A�/�T��7l��}�_�GD?^��c����%�،�b����s�%+�e�}�`Z��U�i��~2vхDu�v����BiB6غa�!�.ʴq��H.����䟛�ᤖ�Ds@սj�k�	������}˼�T^���+ ������E��x�E��;��[BI�1��6�����ͧ�aB�A�;��T/�STg6��/"��$s��}�#ҥbk����݈��\�o@)��Q�+�=��m��g��7�<�<m�N�	�~�YlT�)ܪq*��p�X�;"L���6�]�CéŽ��*/���RlR��H1�v����4��D{hᤎ���/�*(��>��Չ�D!Ò�y�,��-$p��fG ����޻7��ИC�k���F�0�1&��X9��РD'm����-5Pu��m	������([0�	4!�:4�w��pa�T�v�:�\�s�C�i��O*t�!И�(�y?��WX��g�1c�w�wV�_�j<���/���"TQ��E=`�t7��l<Z%�I*�;-��H������	���1�a@*@CD;�<#�)؇M,������?�s��@���i�>~��T0K����*o��߈3f��Pﳶ�ã[tϏ���q�Sj�|ҿ�?.9t��0�[�������$^h�32�gk ($�����` UhZ{�C)\O�p�] fT�T���I���6#�+�q���Ů�t�j�e_�!f+D��y����P$���Vs  &&��ϴ��ֵ*2��G�0�e\X0<��l��IP�#�Lp�T��=�,�
��7M9c[c�6�+ &�,�B���F���[:�
+7`�gA��k"�
P�#CI��#A�I�%4��`�q��Y�����2 $��7oq�4��93S1%Ch����&)oG�a�R�X��=�g�9l$ґ�z�_m�m3jA�����dH���$�����J�*�����jc�b�5n��x����	(��0
�ڨ�!�mHWlz�M�d����ca���rٮ���
A�1`JY���6�[�\G�H���3����G���"k��[L8kDp��8�ZE��*!�:L�Q����sgIW���ƉϬBMۤ[pڻ%)z���j���n��.�\K.&$N��C�>�$65ZQd�i�Zxם� D����NōtE�!d�����#�/�d�0�·,r��4��`e0����>!X��/9�>���6��Vz��@2Ĥ���)�	���.8��BQ��V�Yt�Ӭ瑆Tٝ�*�B.����Jd���!�I����Va��cL��i�J�(��4}�\8ai ���BϿ������)�i#)�5�pba���P ��BE����NGO-��������`�/��x�=��"]��W�7�q g��5o����x=<��z�)%�O.�O�S��?�#�����=?�ǶW��M꿑۾�>�"N_�K��>�����s՟_���K�1���s�5��og>����-�T(*��0�S�g��ָ���.��T�if��'
�B�'rKnY
���k���5��;krTFו���ֺ*Z)�-�F5!Rh�d���F�AEAFޭ�!��$/c�?/������_������{�3���C�|~Kk���?�o��i��i�����x/����x��Py/���?��s�o�� ;����9'������ƬS�e�F�8(=�D�	�*R�I&���hڴYA)AC bZEhAR� �(��T�QJ�5��bj���!=�V����nH�P�P� ���Q�%	HRT�|�������>_���������ާ��9���~���>׆�o���} =_��^��<���/��ֳ���u=�G��q�)����G��L$�;� H�變sZ�UV	H�(� �yH��,Y���m����vs-u�k(�
�y�@��oJǻx��)~�̋���v�ߎ��������q61�ۭ��~621��]��R���� ����ww  s�1ߗ ��g���ĢU��=�e�"[�M�3�5�u�ȕ�&��2��!�h؇��I1�G֣I!�7c�L�i�4.��;�B�YM����O�{�5��a;��.���c�J�
���ײ�6{�Z�N��[�WYSi�X-e��VE�pA��7��ΨL8����"2��څp�9*S&]���0r�9�,N4�� `��Q@-WF�9ٛY7e����ϙ����q{��%SU�#R��s��!&x֞�Mԛ/>]奢�ޱ�B%c_3��*V��amF(7��'���u=G!���䡳����H9�QZۆ�[16z`�Ͽ�ʮڪp��(X%/y��̄��Yr�UV66�X!i_"� ��Q;�VJ��F���N��9\9kk�g%*׭u6(��]�=����2{ҕv�B���� �a#�%T��g͖S@�G� �,�3�t3�}v��D��$����	7�c2��A�`���� ޣR�Џ3�oshh<��ky��2��7��]>���,�o�l`le�٤��e��:������Wl�G�.n3ӝ�2�]@�Ex�Ԃí�A"P��勞9�txƶ�ֱ#/�hlЌɵ��S���N�t�>�|J^�.����+�!�x��ޑ�Z�bf�õСSrSa����IJ��;b�H��N%o�5>� �}G)�clVk���y���6*�,��U�ֶ�=hۣh�]�_s$ �K��t��.�!�}����]ș�tq�ܮ�K�ƒ�Om8�{�ޖ,Ŋ�TI��?z@Ջ��|Jd,B���?6q[cTt�.��m����\�jlH�ƣ��i�ۊ]0��S>ۤ�u��R��@l�l--������c��t4��On0�TR��|GQ�0�5A��"5�� �?�|�&�B���\REyl*��,XE���A��\�m�2N����f]*Nf�΢�JD����H���ے�>���*��R��r&j2t�_^�vD9�r��2P�>FY�M\�-��~hfar^γF �G���m+3I�g�yg�Y��RF��3��d�p�	_gz��)��71���R2����>
;[��':9��E���ӷ(�p�yՙ�ô�`{�k��o*�6=kd�rTt�����`�rN�I,皚�Mֈ��1�X�I<D���N��$a�����$#�#zl�փc�2���_�����d��x7��<�9t���}%y3	��)�'ٵ��Lk:���Q|UO��fJt����ُdNެ����?�Y����r��\C���ş	��Dj���s�����&�Y�f�p݉�CQhJ�V���o�%�7C��냍5�p-�vM��� ���b*�#�>+ν�Mf�Y"xO`e��\�>Y�D�|͕$  ��2�ұ��_������V������dX8
x$(�O�=���}9F �A�"�R!�	�)�s} ��Q<O0O�9.}�-}(㎨��-p	���8Xv��m%A5�~M&�1�X�V�f����EXF��:O�*"��3��U�,�(D�HK]6C�,2�$�`�@�w٦��WJC�� �`&���W�D��b�f9���,��.4�*a����S��d��{9�l,ݚ� yC�x�H�;�gT˸B1�#>�Jtk2�+�MDg&�����
&�\P0�#�"��$BI��Ԕ�
\�1��i G�0��6h+��x���Uͻ� nb)SDK8���`֑@�m7� �e�'+�|���`$�N���Ungi'�	F΋70:�칢.Y=0��|� dY0�x��h���,�$(�(�����r��U��]V.����+o��G ��@R�ˀA� ��)p��=!�� ���ӳ,!Ž�LA�-�S�"�56��#��3Ix��`<a�=��i《#��a8��	jW�(�Vg�T����#1Ȃ���@�(�R��nB����a�\�sB��4��R,ń6��p8$�by)��ъ���)R��*�ْŔ��Id���Z���%8EFPtԅ�.��`u�R�9<�!���v���У��fB�D�$�a� �kN*r��6��>��+�	�:pđ��Av�EG-4�=B�*�$M���S�(��p!��R�P�F��i�,��^e�*dt��Dzv��2l��H �(B�F澵��ĸ�}Q�V�-k���`�d>�������'%`��*+	����g��-�Q�U9�av� #
 M�SKh+�Z�t�������їwsk�_nQZ�R�F����L��,mb�X�"�cDb+DV�lTR$H4e8����P4����/��c/�� #���� pw3�������oس��+�z?�_�b�ֻ������o��?#�]{��w�'\B���9�U�0d �H@�@�2�D�P �U1*��$�
b�2 �TT�bDE1
 h����)B����	
B� �������~����"oa�x^����G�=�~�%���+�[o�w�yGkc��>��:�>H{�����}���ǃR��0�x(Ia ?p;���� p;���A^�pP�cO]~�e����J�-!��\'��"�N�]�jo���Y:º��T��^ ��)�A$�%M�N��x
斺��^q���=�����/i�q��@�%�O�+J��?�   wp�pr� �$��>o�v�:�w���.s�r}���;���[|�:�{X����Q�kٍ��۰�(�;���\wU��pvS1;]�-\��)4ȝ(���|�u2�<.>�\BJd�{-�st>�;&��y��{j1���3Xm@;;č�ޜ�f����GN�GwB!ݪ��LJ]	t� l���u �ctS\CZ�Wlp�2-��Ba�M�MfJcR�(ح���!�>���L���/��)^i]�V��yq�'{��Z޶J#ǈ!��w7�J�\5+�ǃMy�B%ς�����Qy��h��	g"8��v�� �2fC�{#y�6�Js2�\k��΂��U��B�Ǿ7��ӹ��$��0�Ϝ���s�&��B��N�.��3Y�,�C�]��i��*	��
� {���s�SGZ�i	��}���!Z�j��&���t�`$$C�#q���iH�=;p^����f=@�����E�3�_i���H�C�1sBe��px�����±�"�!�[m�f���AT�Ug�ܜ�Ì=Ñ������^g��(ӨD�n�a��X���oR���~�	��.;uܼwǥ���e���^x-V(٨U������r\:M((�����kv�¸r�k�uf
��pJU0�������"�^;ys�	H��X��Q�<�k�9�����h7=s�Ļ��%K��]�)79R0�M�8v�-�����q.*u���
�V<��9v��bI����h���:`�a ��i�$LLO4P�+��`i���WA`v�x���4AU�w����:Jî��>v��Հ�T��e\��28��5M���.��82yq�!��n���D[h�7�'��}褫�n��놜P�b3��[v������<�Հ��}@�܍��GC M��lOY�-�7�cp8Ӫ'3�&S�=d�{��n,���ӭ;���i��}��mqAan	�X�@��s��q- �<���;>_l�D
�V��C�g��m��喺*nqTM�S!�b�|L�%��U�G�K[ڀuc�Ƣ�Z+Fxo/�R��g���f��D�Ϫ2(*�3Wi��r(�˄FK���?�'�>��y���n��d*"�z贵���6.�8F54�B��kym!��ǀ����m� �%�E
�-��ysP*�7Qr���I����ng_��4Уv�u6��f��~0�:_�b��n�0p,NO4Dd���e��fz�"'U�M[�=՗Juي26��B�8w! ,�n����JG����7)fs��q��T%���C����ӥ�\ ����0A��S}�"�$}w�"��ͮП�o!���׿X��H��kP?���l����ѻr�yd����Y���χVu�Z)Yv��%������ݪ�{���b��xz�?�V�7y���p6s�����|_{��y��X@B�!HVS�;7��������i�;5��z�����f�k�た����>K��<�=��i�k��s����ރN{�~�[H��쫠�9츄>�(3Y���:�i�����R���	��a^ ����&�����(Ys�62_vc�D!�E�D- s1�Q��#!	FJ#�o����M�Q�
}�E ��Mzn�ul}-F �6%+�A����Ò>����-�ħ4��t����d�#��Π9��N�Z��%TL���q�*��;g,���*���r�+ H� �;%��`��I�37�(�Z'�����������V�
l�Ӛ�D�k��6�Yd/|ͪsN ��8I,��E����΀�Ĉ"�*3��P�zWG��`�:hT%�o �0G�@`IlֹeS��-��2ifBqf�I ���9-�U)l0<�h�2�.Z�2j� Q�$撘��Fa�P�j6�
c̯qk)p,�'�h�-IHI"�H~��D�n"��T
 @-x�mAZ$�s�pƤJp&c+�ke
]0��Gb��T+�8�B�o����`q>�'z�G�:���G�@p�Q}�M#��]����&
k��z���ഖ	j�b��6#�XP����@$L6ǘ"+��(�%5�Yp��U1�\.��VQm�L��aOuQ�(�4��Î(ҏP�A`�	S�"B�8�0�V�iP��|�<�(@aS95��y̥�A9 ��^K*H�������J���XɃ�"Lz��\��z�\Z��'Fph���p@p4�J�`:�lN	�Ǩ�# ��z���.d4��
A�q4	h�ۻ�j�E�M�h�Z��j��xֹX��EsZ�ۦ#BZ5�[�xۦ�ّ]�Ѵn�M������t���~�o��:#�}�%����ߺ?�����?��m�~g����׼�o켗������^��7�x^����O���������9��ݸ�'M�}�����^����	���5�q���v�4�h@6_��^K����h��+�{Myw��8}�}�}w�/�-*z�}�${4�g���+�!���})�s�%�������B>��^�w��Di����W�˻��	���-E�ZG� �$]'��ު�/�P��m'i���n���0"��1��}��� �{��Pq��ᆹ��ne�u�\�;QWLu�Gk��+-Gxl��Er�<5bp�����4!Y�  ����Q�;{7t�t��(�����nP�g�Bݚ����܂�(�5�b�$�/s�X���7��oܾ��Ƿ�����$�v����^�b3�fu3|+n�j��tL���i<�}Vƛ�ig������*Oa2��!�9�w��M��Zo8MX�>z�?�@��Y+����9I����-�>xE�e���V���e�3�Ι4/,���j>����L�D\M�$l
����H@b��Y�P�t�_@\�F6Q�0��NS�R뫶����%/Ik������00�-M�c�
�F��I��(���fI̫rn�u]�{`^��>�SnGG�X�0�>h#^T�.�T�@�t�ʒ�a|p��B-xd��N���w�����M��?=�(�P�����.�c	��I	�������w��K���`�c�U��|�ZD�+�]�1�
��x�����V'-��p����|�^N�;��?U	P.�5Z��5���⑕l5�b왶(u	 ��QU��#kbt&Ad9���������	�9ɪ������;��$K�Eq�4�O��L�]��Y,;\y���}оb
�A�8<*�&+��k��/��Jm%�N�}����']����d�Yў-]zF���� �ݪD�`�t	6�G+�烵�E��d�Qe�{��_ە��I�$B���+�&����ۨ�Y��^gL����ċ�����������#�I�F�J��F9�o�b��ǡ���J���l)�+�۩g��2b%�@�ݠ<�l�) Hjrz`�2g5iQ>���[W������[JA'6,��?���qeN�ۻ>�j���9ѷF����Q�~�onf3@��E��Q�\f5�������a�>�wI4��۸MV�v?�zè��^��f磖#$�Eq�w`Ԡ`���/s��o-zw�Cdp���/��[�j4q 顣:A�aPҨ[��$e��	��jq:tl�eX�-����J�tq���᳃���P"��ʲ���7Oy�������*L�ES[��r�)ǖ-�a�L�mH�n��u�q*c��ƛ��t�ce#]��Hx��O�����3B�4��R��/\O<���|�,핚��h���	�H�Օ?�CH[�͙#�7$�eP^MlBM[d�T���"=M2�����>�1q;�X݀�L�I��M:���V�
:���[���8����B�𳣖g0Ij`xԋ*�N�%�)�r�N����
��jo���7�_kL��%Y��5��)HN�\�)� �j��ŷ>�	���q��d���AȲc�8�A~7A�.��n���g(i�5Q{�M�P�EY�Ӽ���q&w+^�L�"�f6�&k���2.DG����0қ���w��>,#��q{�����ա��߉�x�M�yOu����O�~�ڥ�� b|qߜ����	Fx3]prL�Ҟ{%['V_����Ǌ'�v���.��?`���,LC	�">����/<�� s�$9�9/�|X�zq������{y�.:|��X��k�_i�jN��P�R����>~~��aFjf@�.xf��CL�Ʌ���P�ʁ���:�IN�	dW�R� V�S�2i�jE�$$��Uk*s���hI:(L�äz�j�H��m�N%�PEd(��-�L��q!3F��8�j��Ð�D���'7 ���N �D	�J��Eh$�+Y��@�h�Fq&:�,	�Z�.p�V9����+����TV�SNX�$�[!�Z��%q&s���U��cA�y�>��9�>�f���'����g�y���1� �n%�$�$$�Ѭ� Ɣ�2��M<�� ��
�qQ�v
jp��A����R��J\HV)�f�M*.
\��Ey�RP�ơ@u�E5H
��#R�z<%�-�hV���[bM���%�����O��R�j�����l��l��|��:v�1ɀyt�����0����Ir�J�Ƥ����T���4�2�4a�a_"&�4��A����e�z�U"�VC==S��T?/��>�w�����*���9�Δ��^8�\��������g��󝣶_a�\��s��>��  ``0�O� ��:�J!���,�v��E���'�\�v���]��`��L�ۺ�J�+���mtl���sh�Tj
ŋcRQ���/)E�̓��N!+IGO�W���o��杚���aW��߿�?����������[���\���O�����_[�������\�'�����7���N��?��	&���nc��Ǹ�r�l͗&f��`��$c�ѳ�n����p���Ƙ�j
q7��ooE[���b2eQ������pcs����QÖnsk�64�\{�f9y���xh,����q�o��}�vA���$C�ݽ[�^��\5���3B�Au�ܯ��Ul�u��V�{���޵Ov=�w��r�|��B3�<�pA���Ӻ�������	tS��t1ݱ���dD=.�S�.ۨ�s�l�/[��L�_뒡խe��4�隖��̊���e��j��%t�]!�դ��Mgz�w$��%um�� �>+��]�ZwH1p:|���T
�Q��q���2��8ܹ3$�uw�Z�,���c��.�;��̫�9D�v���������y6�̜N������:�vɚ��Wh�Q���n���&9�6.E�+�X������&<��&� <>*H�|����Ǚ�������^��{_��>7{��Kƞ#��7��GW��u>�������E�B�����/hǺC�C�E<.����B�O&a�n}��2]��B�	���'���ѱ�g�o����Ci5E|E��Z����C����r��J k�����1���7zZ{2n,j�/e���)({�%���������A������MV:2�����܏.���"!6��e������w�G����[���k1w�du�]=*X�.���Q&P��Y�Z���é�8��u:�L�^�j�\�zExQ	DJ`���k���w���7"�J��G�pڷvG�t!��}�h��N�p���*	a�f�8�M,,�νBxt�GV.����B�6�tj�6bƥ���]9�'2��T.�N�aܻwԷ3/1Z5ü�^��س� [O9�\)+������lt�0��ٯ�(�V�� �8��jd��yo�gN�?��dZ#l��\�
`X�Q����.-\
��A��qrm_V����n`��-"Τ�{<ǭM�5(�ö|�T]���ő�:�.k�jG��ə�WϷ>c�BM��5��`]V�d���-̈́�v���1&	�� m_}�0(Q6X�4��:F���۷����>a@��k	T�ǟ@�ʝ{�7>�w�	GLξ=Pv��u�2���.�#z���,E�1rf�_���i���_��u�����H��NM�bd|w%(��I�1����j�)�4����b�H��*��M��Ӌ����V��M!
�h��ZK{gDal��!��������^�\X��M"�u��CV7 �m`CJ�=����m,���(�>Z�ΖW��v;r=4���+�m��A����=%����R�iד���
����BA�p�V���M�����8l؝*�r�J��Cpa�k,ܞ)Yβ���:[7EÁ�d���d|Nwׄ9w�A"~B��ld�@�J�����e�{\�1�������o?4�d>sj|��|�o��s��o��� 62(j'��	+c9=���c\�k�0%�y���	u�Ƌ\���K�b�F��-��u� 7�Q��nV�U{}��گ3K���Gcd�2�̑{;�Qa���汱7><���U�"gp���F#ˬ�՝�w��`�p�n*�\��˫�.@~�B������c ��*A{�2�z(��v|�؟WA�5�H���Fܛ���Ҟ<[M�Oj��ilj�����$Z,����س��Q7��Xڃ�����N����!��P�]�J�^�NK3yq�|����!��[˄�p4ن��:Ł��;s��5��J��.6kv�Q� ��D,;P:-�������e�� <�j'#fF�S�@ժ��÷ML^5�|q%���0�m��`M��He'���$����v�A$X�`��(:��msxz�����g��&������xZ�ݩ�t�U��\7eʼ���Z�FB�v��i���T���?��l�ajo��A8�+2��K��(K��[����J�!�[�hu0Cl\,��Qs��n�G��a �y{;1�6�s�De��T 1�P�&���#v�^���^}.׋��̻^M�1��LJۧp��y����G/���{@�7�1 c�}���aL�|�h1DĖ��Q��O��~���<Os��
��~!���M?,Z]tK;��}>��=�c���M��:{��t���p�(���Ov����U�I{K㗜���1�_�Ն�����!yK``&C��$̛�ꪴφ��Z)H��N����:B"#8@
2jL�"�s����2H�̏���d� �鼼������	���� ��	6��\��2%9BS�����喾�;�?0�|�ߒdZ3��&��::i^���S��2�K�A!�I%NQr�8� ψ�%��M��Fo�j�~+�*�s�sOS����T��|a�������I.�/ϕ肋%j'_���Q�[Y�ϓqh��^Sq�f��z�_ǧ��?�|�����������o\����Q�}�.��秾�)��MeəsG�RJ!FhVL!$S"�"�$�f�3�,�b��h�ɩ9��Q�5���Nk��g�-��|"�+�7�U��i���U�;)��oٮ�([{�ze���?9��ҿ,;�}����y��hV#�t'2�HbA-&��	,)@ԭ�QA�<��LM>�q�[��V��}>ۯ��+��s�����g�$,ǰʢ��<�<��T��!IEKcI�*����.m�ͱ�V�mͭ�\�se��nWb,5��%b 8x0
�>�p��=��>�a�>�~)��Oo��������:��~?S��~�>���/��:�����k�{�s��^��~�����h �t�.����ݼN��7�	A<Ȥd� �0�y�q=ۄpq�q]�S�goAqۜ�܍��]R�g.�`W�62nÏҮ��[���z����/�lR�Њ���Ќ�Q�n�f�F������Ի�59Dd�Y���N[Z0C�����axk�۔����՗p̫���/���,����{�«��pL�)ڄP;U1w���wuQ�`�7�P�y��3�2�d�enfI�p�]��uv���v+���%���cd��!Or�DT��ys1-�O��L�p*�.��zL�_I��p��s�-��H�nEJ��G��)!�F��]�����o{r�g+'���s.;�w�,'m�_���0�u.v�I��y�����n[��Y�7v�͸s�c�Q�y���VU�g`�-A�:Y	l�. �ŕֱc�lU�\T�s�=��r���.�(��u�(GS9�ڇV#a��dZܮ�I�߮��oD��|��
\��S�`��/יѪR��D��:�T��������ѹK���_/hi�ӽ-����ګl�ą"i�vUD���(�X�R�ۋ3y:S��)��ƻ&��Tt��*��l��YF2rs���U�y�姵�&�sݕ7l��ܝ�0c}�@� ׾��+������
f���D�]R3i](3�7�j���\NX�@��w�g#�f��q�l �c^B��C�/W�~����d7����=7�{M��������z��ޱ������;����>"ǝ���~�&��(�u�>l�C]�<��z/%�=�sx	�(%���i��� )VhF��!�������T��h�A, �����������)����/�{��d{��<DV�3�Q�&��<h�H����"�?7n5����� ���޼�B���4��~�=5]�ÿ������ج�EVɰ���-��nʫ[5���/:ޫ�n``���0�k �~H
�.�.�'�B��8��K��#�^:���#O�k"x��nV�N��
�:�`�y��>�%p���� ;7��~E��B�g.k�/b\^c$�0��S�[ @��ytZ��eB_{.v6�$NV�8�6��>��#��U���K	�l�L��uj��P3	�P��3�m�)>����>�,��'�'/���&��ό��heӏ���U�Z:8���
��e�"�J�s�'�s�Uv��sE���A.�z��t��q�KS6u������xio�G�6p��r�����۹��~wu���0�x�F��E��5�S�B����)|�����d��r��d�d�'�t+��?X�t�O�:1�C��������&]�������~�5W��w�b�L�9e#q\;C$���P�� ���72�~�{ f`[�_��2�G@�-?Q5H�{�Y���m�L�q�n���!ݲS �;x�_B�v�v^O�~�Cy�������A���QD�����p]VM�hE �uN۩���d����8��E�z�*6��ݖ�lJG)حx��'Jx�F�F
r�X�dp��dB�YtG͢ndՂ�W�.�m�3�Q�'�~,��qNÎ:�Ѹ��7:"*D��3�%	�T�-Z%6��o��G"���J�P�Ƿ6,�Q'8��!=OǊ���<h��/t����r_�O�!�J�����%�$F�C�xL��\Ͷ�ԫ�(ld�gs�k9_|�w~��auVYA�cXs�R�ə#�͕�Ap�g���!�,��@�M��"m6˯#���I:�N�$V��+�\��tƙ�2�颣e���D4.f���q�.���5�����,X4娚&n��XuZ8j\m't���M�hWo1�&��hYR�w ��u4��MQ��t4_zC$hP�9i�)`���fA���x��(�A)��J������ڜ��~�_���>2���Z��,��٤܎��_6��)
�oM%sx�+��v!]I�n)a�留�;xs����9���7絵y�����g2�=��W�h�C���Jf���U{-u�*���No�Bݹ
W��֩��8U]���QQ����nZ'xɯ�.�]U��R�^*X�H���xO�D�x7:7i��ip�%��Í,����S�{]��U 9���c(\F�M&��̨�Ch�� ���:�'3;���5x����5�+��W/��Ӹ�wo&]�ȭ�)Ytٚ)�E�GOqL�Uo
�Z�W��N�©��<dϨ����wo����8������PH�U�
��/�Y6��f�f�_��r�  wwb��0XB��@0�h�x�Vo-�����}������;�	S�)��N�� �#�����w$j���S����(?�k�����+I{��Hy�L�ҥ�ߛ��*fm�ܳ�ƴ��������^Η��x��o.m�Z'|�
�ZCgV���������U��N�z��/=���/�4n^��輕1�+��Y^�������m���&]])Nʋ��pN�<�ܯ_7|��g��ozk�KL�Oyvl���n��˾^�=�^�=����z��-J�-�����N(��;�/�Ϟ��{z�
;w��'
)��Wi�8{N����u�;z٦[�궕L���=ݷ?n���}��u�]ĝ�/Gp���,Xr�s������9{gR֗��1E.|PI��}}}|_Hl���>��{:=���2�׏xy�����Oj���9��_I���"��}}k�î\��6�M�}9隧.3�On)Wڡ�AM��k-��)r�}<�G�U�$a���-}�����x[���{��w�nO�{q�t�'�n+/]ۼ[Zu��_��o�/8�˧_z�v������@?��~O� ��,�c��8a��NPErU:��[b�W����ZVW#O�jfƱjME��nk��m�ռ��wC��LX)�<|p�F�^�����՗S�>7��܇������^w�9M]Ga�������}�����Ϣ��[�����m�������>mC���@9�������#"ń�݇<��80M�a���n��l���3&2�1AL�F��cS&L�%�Bd�(��!J�����^��y�����B��@+@� R! J9�|�}�g�e�{�V�7o���O��=O��>{��p���t?��O ������x��>�h���< �G��|3��J���H�G��=ç�)F�Jo����g��2�w>���� {w�%C�h���)�El�����l��4����o�ވ�xZ�x@��9���	��.%�̦H��ȓ��t\�KE��uly���X9)U2;�	�Xos�����9�����wwp]�� ]�p@ �#�b0���H}�0��<cS��]���B��iͷ�9�=�с����C7�gJ���^�_��Xh��;���3��]��V����5-��Y+W��T��"p��Ç(��v���	��:2Z�b˗:��Уܙ�!�JC�)f�L�,��[����R��ݑ�xZ3��t�l�
��,�ډ]�e`§Kf͋p�$F�9��u������h�ie��VZ�jQ��\�䰢��'�ޕ�Z����?4ZH�GWAnR�^�n�����7#q����S����'f�exyI�m���Xxm��^�I���n;D�am����شP�7�)�������=춧\c�=bU�ּ�2�z��
:
n�0���f����N�뷈j`��u�O���W&�z��V�94}vh`85>9����	3?�����ھ�J%�Flȫr�����t��Z;g���2z�盳��� <�����@��lܭt^t�L�7���&ry)+TR~,�qY��$"1�EJ����n|ZxJ
a�΅��:teή������|�%պ��%!��P�s�c��2`��p��"N��Qe�������H�D��H8c),�|�ݲ�cr'����)+[�`���>�)�q����&kE
�r���0R�l�SD=��FD��;t���s��`��ڐwP���t䙒Fn����'���e>�o;jWƱ��^nt��,ʴg`8�߂��
rKA�FX�Ҧ(8&��)1�Zku6�i�N�|w��z=��-B!Y҈`�)ps�~���
"xU�ʜ`�yCd��1	���K��f1R��OJ�(�N|�aQ�p۹ź��bp�Y4�jf��L׋�Oc̨��?�	��'���W�y9f"o��ꗋ�Lg'�a�^�\�'�<����N���j\�s��C�����3��|�p,Đd�QJ��bTO�?�:��k�Y�U��D�1t��t1��n��F�>�gg���7��2rxl�a�a(��wsۋ�c�Jm~��8���Ŭf��8�!�!.���6h۝�0�I#0su'�w0(D�h��
]�tOX:.ʆа���������;�T�{w��s��FSt�~Y�e�ʵpۚ_%������8��{������J�`b&u�bd���a�l��nM��Tqo����{��˘Y�m"��m�x�� ��0 tT�t���T��T`����i>�V���.�ib���;t`��+o�
�R�1	��BJ���,W��[���dK|[��J\�B�"n�&�����	�g7XN��=a�3iF=y���nO%���4Kb�D�o>r#0�h�nUc�
�i��;�J�?D p;�w�.� ҅ �Py7�|����[��|�9�mi��v�^٧�g��x!��A�>��
_q�?�$�}���%��=��x	��=����&�2/��d[^�W����:����B�O#ü��M�I4�:��ͨ��tT�s�/��[��S�pw�2ϗ\������x��G��5���{N��\ۍo��6����y�kaݺk�Zp��:�|t)˾�?��~)���I>�y���^�>S�t��x�n�SP�P��o�֫|j�Μ������祼c��Xxk_ˣk���eR>4�_;t�w{�5�o*�[�i�5��>z�m߷xD�x���PYL�{qE�qM*,�!:ԮG�8~O�k�{k�ow(�~����+wW�{O,�~+�,���.�m2w[9uʡ�/r�l�]&!)(�-�',�>���̺v�v��Ѽ�Uh�}���安H:/\�ݣ�U߯Z�~��ݼ_��Ɂ��` ?�?� �$���F!O�:�7V"X�����E֬�l�o͕�Z6�mDm�u�Ԥ�*����X�(s����-_���t���x������q��s��/��u���{��t�/�𼿻��?��zs���x������1������;����[g���C�t6,D����7��%O�����&TgFU�X�"����Qeؾ��w5RW5Qr�%=�o޾��=��Մ�����
_ش�]Ea<���[�f��E���j�pF���7��E\.�6�\�f���X7���d��ˋ���к�9ok�ɽ�#��0a�9�������T[����땋���."��enlr�b�Ek��:�Ć��U�ۚ�������>�XΫ��_��ܳ8o�7`N���/�D���di��n�zu��w�:໌�spƩ�'h�1\!��^9ުI(<uN�G���U&�����U��M�rh(�]6��U�mͫ�~NI��-�V-�yRz`��O\��AQsYy����\eI�����ˣ=d�Q
Uc�Wfci�T.���N��j)YG�cb�s}^�z�L
וFx���{��QWw�J�y�܌H�n��b+#yͨ�N���VBffʛ�^ͦ�؜��w�^-u�띾��gU�|�ϵ=��Tt�9��S��+����{4��m���yp	�a�]i홅��ż�[F��#9��#cB�{,�h"m��6�n������Ι�Z�����9�y�q;�ʇ3��^en�Iއ�&�#����2��4�ҭ�ó����Ɣ��´���2js��eb��6�1>v���Ȯ�V��O>�jɶ�y��_}��Z%�Ou�T�Ju`�w��S��YP��03{�z�`�m�-�����]�%�����}��J}ֈ�ѷ[f�Y-Ne�ꁳμ]]B�E�x\	{׻�t��[�w1$s-��'Cu$�,�lp�j��C�����yr�xj\���n-��.L>e ٸ���w�-Og���7gs�#΃|/���Nɱ��jj`��de�7���u��1y��1���hҡc2q8�&:'�kF�ԯ6ɚ��-��MiN'hFf�A$�*d���E{5��ٌ;~�LF�FYY ���ˣ[{��	��؞ws;t��X:��\$�FEn�l��ݼ��8�׍GN��l��с̩�k/����Z���������ϠFL��yWѩ�������<�7������վZ�\�)�qۙ�13v�J&�4psZ6w�����c�l�F���<P8˝��'GX��d�C��I�2/'I��1�S
ȩ}����;��\�"��><bؕ���Ҝ��}�0�f
���t���F۸�p;�.�h-չ7YƧڧF��yu����;3��]jo�½ڥ�ؼ	�_t�^�l˶�n"�A4/=��Y��;/�m76�B!R���f�g9�=v�fZ�ډ�9��a�͊�6opǛ�#T����F��t���ם�� �{�dvwV+u����7�y1��_+�{*:����g��ыt̚�]v����Z�ם�[�"���e�V��qGB8�;�gf�.w�b����"�e�YōȪ3u\�]��wQ��
�_�VWVnہ�w�;Db�D]D���'>���v!���M�����)Hձ�w����sA�D���ٹ�ƺ'P�P��L-Ȍ����r��0����o%��٭���V7r;9��:�M^9��C�ݛs��d�3elN�s| 0K&b�bXb�B��Sl̪���f���r.��!x��2d���sx�ܘc}�awiO��o�b^7s5fa{T0=ɮ��po'd��̈́hh�B&��w�V�,�4�@71�{�[;�\r����x�g]u����k5=޹��z`ݦ#Dj	�x�̑��U33w�#N�.��?"\�����mΈ��Ss��^8�[>�$VUáч:��u0��=5��p`N��k�\���������՛��Y��P�(H{3J��iM�V�;�'k;b�6f�],Bî� ��ѹw�t�)È\��*�+�6f(�w�w_Y����gL��
؎�1�����S3&6�y������]Ѫ���͍S�Q�9m�ܛ�CӸ���dV��>��U��`�G+�m�V�곜�!)"�]j�oj���iF��7���-�=UԘP#VF���^Iɺͪ�yӢ����F��
�3b�gTugb�g�nDm��u�2�v�h���,���0`L6�/*6kR�M7���.�b&���Oyw���f�2',��b$�Ò7j�r�{�I1�ú���:��nJ˛��]��G��]�ܻ9ǩeg,5;aS\�^N	SHtP�B�\ƅ�w�s��`��������-�X�q���Gh[��8d�;��qt�&#v�VMs���
�;f���E��ᵛ�&Kڧov"0!�n�[r��8T]
ٜ��w�L)��o3�B�p��u�(5�/�\�jqk͡�yc}Fv!��nQ��TG�z�D­�D@�[q.Yq�:c��T@g�����k��gÄ��Gne�O�EZ��Ǳf*/gna]d�u����[U��pV��0�y�l�'z6�Tv�̕�QeJڜ��(��TFn�(�C{R�w��q�2�8�A�����"�"�����[��3k�7��۱`�+�j���6)e�.�%��lp����)�Z+�rn�ehz::�؎�.�U=2�����lon�򝮜�x/��5�1<�f�*�J���,���\�\C�ת�@�v��ŷ]yW�ޫ�y%l�t���fU�	��pwXו"����Ŵ�-��U�ѦSƷs3���9�pW8rҪ��;���+��r3B�1�Ċ���ڍu/�"CM�י$Z���,��s�Tf�V����4�l^p��}�уX;j�i��;pc�"q_8�1V�����&�K�f�z���ڇ�Dt�
.a��[a����n6kfa��.�/�\..����`N���<�[���w>��k��>�d6�	�J5]���,�]n��Ub�T�Q}��0n$�gf�\����o*i��]���ڽ�y������h{���{댧uc��fU�.�jƍ�=�V4���5en���FTL7�)f�b�h��Z,�[л.�l!x�hfWc[0��'v�no���n'��ښ�XC�=�f�L�M����mr�,mMѭ'Q�l��ܦb��t���
�1���W"�S�͔��]��giF9�A]�b]�,źf=�z����.��B�!V����4*������r����뛬�Nw�ik,��w�wVlȢ�gh��uܝ�M�����2)P�,Տ{}z��$wC��렒̓���q̚�fO)�M��q�:�=FG��%���aZ�����Éo'�\���=b�0:x��iw\��\L!�2s*B<7�5e58:.���x(�^9/���	o=*'�ۻ������c�\�q��c}�jC�S��L�d��DE�1�\;�F,A��.�Tn%s[�mqd�C��{|o�T��X"���$^�f��s�)^CRs%>������3�	����|�5T8em=�'U�����`��ֳ5�c/��z"!=����jvvhlDV4.r��U�U�2c*D�w��M���{\��c;.!�pUw=�C�XjVgao������wj��59��̤)��lE�zY�p���]nݒ5��lt�k��Ҩmc��۾"�9F����LG�.���,�ە�FA�;�=��5�u���j��f���|ϜM��{-\�r{�]�q3|^ N�P��Xrʮ�+�jk h��JEIjy�+%,]7ELm�<��K��mҙ���f2t�]��;����Wo$���@P���a���4�.6�`qϓ���t)���(.��(j�UM�:8Nf���]�v>��tek���_���n��ޭUڌ����:%a��3jS�3T5�G�V�{3�Y��Ў�T���Ж�T��2^ʎ����1���a��Ӹ���t�[��݊ћ�S!r�5��GN�0�,h(�љ˻D����;�E��˝95B�����y3%�ws5�������_��W�"�=�˶�V�х\���n���:��|l�ۗݢp��`�ם]::�Nͼf������리N<����d�u�b��}���-�Q;��j���XV���n���	��d]l��E�%��UEч�DH���\�Q�Qf�a�D��2��."�@t�/ي�Z�|��-��B�I륙�N9�!,��]Gg9m��v+�IU��LMJ굽��������UϓEmmV.�=@��٩1-"�{�������z��&f,�e+��hl���!ۺh�Nf���E�l��w(FWb��q����i����c�����2����u3q�����;Hҡܲ���5v�S���݄g��v6Mr�g�D�L�wr边{S�w`��[�rnv6-��u�4�R����7l�7���q�i꜋����4�;��˞�8�S���.xd��4�I�!񧝌V���b����E��fe�ڻ�@�Zqfc����d���#6�k
�	ͫ�"q�S<n�a�E�v:0�>���K�B�;��a�f^u׭�wA1"6�Lxnt�B��Hů�U:�"���l�B�"�f�=W��9S8y��Ӣ�O9�/f"jY$��*A���U(Z"��3o3�o�K�3R��r����C7#�f�����[�S2��;�(8�Mnl�.�0��Y=ʞFsm�в�+��՜�/�Mi\=^������=����P�=�*�="*N�ٕc};aV�=���K��ۇ���۝�s�.�aЋ%P��������t�W��fj2n��ٽ�bC��d���q��}D�U���4'jiQ�����G0���4����[}��Yu�EeD����^u�h�����պ&j/wR�5f�Ϊ�����2��̺r�P;���%y�CJB�Dp��.�ӶpJT:*����^���UZ�d�м�/7GGG"fuLY7gf\���)s���b���Z˵$�ʖn5��Y:��!�.�da�**V�ڼ�t��u�Ȭ��]*�(���B��D��18��ꜭo7n�sR�=9���\�M�FE��M�����ޘ��5��UU5���t����[���T�SJ��d�����`������Ǜv��
/<8��J����NE�r�w.�`e'SCf���lT���,#��Yxhe�D�䱉j���.�������E�P���c���>��9��FSC<6�<���[l��l9V,=�f��Y\�Ѵ�@���DȹغWU,�7�N]^2��q=��^b�u����u�[Tko���^<�rL�8.��槹NZ ���V8�S�c7:��@�Ph��5y���sV^!o���$�F �(=�LL���cn�[�=;s'C���u���ٍ׏
��M�;�lZov��˳٧������T�u�J��VlT>ɽu�5'q�~1�*����U���tN��]�A�8.s���/^Ɔ�7}ִ�FK���XN��ɩ�0)�/)��t�{�3Eo;]Tg`B���.a�U����5�U��1��۪ڪ�饆rbl�+�,�N��s���������X�+�:�h��d���7F^�1�ಠ����ibN��&Ҩȓ��w[3աl�As�)�+���,�d����T��q@�����^�r��%bv��^�x�]�N�${*�?rx����A����Zlfb��Osjo�R�gT^�;���o]�/]gQ�w��w<.w�`܎Z�����Ե�N�g�,ݍ�+^��ڰH܍U�dIX*�M����6���yK2*ⶹj���
�7g��)�;�j2u\t]����&gܮ����Qٔ�r1�WS$M�t����3+ҹ��F�p���DE�V���b���I�35������2w�ғ`ZP������.r/��,r,�S�mF�by6R���ݖ�D@S�#PN	�Uwۺ;�|�ps�
����p}!�he�T_i����Yb�B�8�c2�é�٘�v*�S��sj�iٚJ���#�'�d��=wek��x�HO�9�~��͈��F>���� 9ӛ��ɢV�X�N�n^s�މ�������C+�kvr����{\���Qڔ�'���8Gjq-��闧"��R�=5��(l��p��
�a��.��:Òř�ʷ6���;z�"Pz�mY�p!x��ٰT���]��Td��̩���d��N"f2eWHՋ�z�V\2e\�Cv�u�D��dm�o��<��;p�)���}��<��#�w�|�(7-)R�}�p����fh�!��
sB*-mZm-��FmX=d�tq�=��[��ަ���ޜ&�bL)MWU[�֑��ຌ��9w��X�����66�P�N�3q���u��n��tMm�®H���6���wYS�Ԧ=n ��V.9W.�D�Ǒ�9����j�ng]ɞ���(ڵ۵#W
�bs��!nH/8;�U_`��V<m�(�\7E�W[�&/���BVm8H���d\eb2&n.�<��[�/rz.�/"iI���b�]�r��;r�o'��}�m��"{+̈���8�ei\�;Ń�u[����0a*kS�$�J7*Ir:��9;�"�訨응�[�Oz���A�8��r�*�d<҆��}9�\{��c*ͣt0�{z��{x���_i�DR�`�u�@�K!���}��Nн���a�H��S��5��q�������47}��8���wv���JqJ�c��:��yɃ����CǺZ��w�oʙD*p�z�3�.�YS2��W^�m�4Q鎈�L�qE S�j�Ǔ���ڍ�I�f�]�������r{��LW�ī����Ƿ`�}3;�&}�J���y��̇�sF�lf��I&'I��ECڸ�:F+2:�bˣt.��Ug|��&��ܡ9&H7#L��ܹ-M@�[��*WW$���u�]W5���gq�p��E�<D�6�o�숊�쩽�+����UZ�;��6$FM�=+��levf�;�s&�gkg+i�/c�>6&\����:!f�s�{w�.2VQ�մ� Y�������['�M赪.#�m�{yr5���*y3F�4�Y웺؀f���Ev�{CY��bf�Oq�l���pO8<�1��&��]7ih����W	��ȳ�,�Xs�-��R�Onm^2�b����lG�Ub�&���j�ވ){Y�d�zk�R��!��s�Fh��gq�F�V�����]��uPz#\ܤ)��U�6o7��FAsy[թ�\�F.��r�.���K������pr���Vrb�h����(��4�)�\H}7'&���v�F���u�u*�5&rC�N�0��1�eI��n�"qnXb�;;L@�hb�*�NE��;��D�WVf(;r�����������v�;�1�;���:2�nf���c���7b7�3p�XA�UQOU\�3q8�i[qQS|҃�OMY�ɷ}��˖hO6���sr�;��Uf/7N�ttlLV^�\�a���V,}w�f	݅z-q���VVI����������������8�/���y�}�\��7��6������1�}�|Y�ōڍ�5��%�d�d��Db��[�Yb�#JA�X��!�A���g%ۑP�&���D�%֮�B�.����Q�f:�G�B:pgh�7Wh��(��#�����tk����B�al*��3�(Ԫ.�]g ����q�7]P�3R�Ѯ����[q*����B�/�һ�{��������wejgT�t̙��GGOlR��V�{�V�:f\�G�jhu2��<vN�U���������/Nr�c���{jcۼM�:�X�c��R���M�ۜJ#Sw+��1��.�V�t�ȅD��I��n��F�T����t�#_k�EfJ8fzka-���=����U�ϓ�H�}YY{
rk�m����(^�.u\yĵ\mC��>�Ã]g���L���2�@���"��3ѝ={�d�B���;o�U�]Է�JlX=�-�s*�ә���l�+�cޘs�8�9j\��>-<�=���UM\�1ɭ�11|�1�!Y���V�Pk1q��ޒl�f���VB�n�I���gn'w
ڎ��&j���b���(m=�b!�(��{���d�����qT��辻�j��-rc%�Vtm�nv�y����/���H�t����Au������NIk�\p�䰃[Z;fg�Y]ugw��̐`E��#��R�+3�hO�v7�̥���=tn:��ͽ1F���[U��D�D�;<vj��nf��;��'_/H��3��;����������
cW^��y���k(����шR'\�POnU��72���<�Q��x��5��Q�r�nY�J�|�Oa�Y�G���Nw�7
��7���մ��]�r���˸�<��ꊌ);���e0�;ga�։���b.D�J�6�滬�^,�N*Eڦ�����L��D_f.D���y
�I�N��b��w.��{��z�^-j_��=�W;B��cPQҎ-�]�yq��8�,��W&�ŞU\���T�}�=�i^�)"�����sڮ�b�0DU�n��'(�M�o:�Ex�l������L]S˲J�.�V%j��c/��!��(m�4��K�U��j>r���w�w/2!�f<�vt���35���Z�g�T3�j�vU�*�����ZgBǮƎ��yS�ugV��Nsz�k�� �d�|#S���◑B��ШVj�������.J\����n�����g��t6���/C�5�G{�E�[�\�_fO^���Pg��������ٙ�ɱ8�����V��S�7�k�[<v_c��]T'������.Iz�"����"z뉚�I���U<���{/��e�Nf�ލ��Y��r�\�U�zp�k+����	�)�5�tv\I�JVg%fܗ�o�v��R,U�D�_u��e��z���z
�ڍNdd��P{��;���"�tu���s�*zWE6Y��\�mF)�$��;�KF��#����3ӻ�\��C�Y�NN�鹑|9M}.	�j8�YU�Y��� ���_v��hV�d�3w��e��@� �� O�y��X��)Ei�B���+wvأmr�kwW9�Qh�-nI���6����6��-i**��Q���LF)6���#�5IX�m�*���sq�clTj�Ŷ+r�����6��QTX�U�ʪLkr�w]��+��TZ�wvѪ9k���Fբ�k�.ss\ۖ�g]��栢771� �E\��.m�sS�F��Qm͹lZ6�ݫ�Esc���s\��r�5Q[��jKlU�m�W*�V-Z*ܮmHZA)�Z�hbGp�"*m�>�L��쌣���i�|�ާ֐G��_H?��=a
k�}����2{�x��ڨ���K�������{BYы����uv؁vZ��{ġ�$����%�+�W�������'Y&��m������1d���/��v��=Nc58Yw�E��%2�����H�����(�����*DjXN�E���n����)Ϗ��ݾ�D�ɏ#6��ЩN���zS�B��Gp ��"�FyL*w���`5���|�j���i)���bV�n��������g~�Ȟ��N��hw�p� �$e@���6�78p�u�gYI�Z#�T4C�)����k�J@�N$^lv���qʴ:;�>C����^j��tn���|2�:�pYy5����k�4��td�>�U3-~^u=�r��bс`܊��?��X�/<�1ډ���(�ƙ18jY��e�)�G�dQ�(�5�,,I^�Q20�ʴ,�N��A��/\�N�Cy)���V4j�˙�:5t�d�.7�ܣu�L�sK3'�n�^RS�܁3Og���SwM�`x������K-��ۡ�[t�	�8����|�n���_����<��l��0[���7|�+M�Od�'X��z��dA�Ij]~�;�GI^:�A��g��v���87��چI$���U�ڷ�W.�M�T�j�'ͅ:K{�Q��o�n�l����=lt�N�2�/l�sx����ō�n<ˌ�K�M�$��WO&�R�9���"�F�̃Ϙ�M���Dws���,�M8$�=87Yu��8��7�N�թ��n 9��EN�����r!���,��o(gd�X�6B�L��:�C~2���L���)����VD��ؼ�!��T��7W+{u(AGzU��k��<��SԊ��P�F���]c��u��^�|5e��	&b�E8'Xݯ�Wi�C�6sOU�w�����4e�\`ϋ��2#t�}ؽ�Tև+u9 ���`kA�;�5�+|#�cN�b�ˏ��P�tdQ�/(�{���(����pO�����H�HL��^���Ğ�br~��w�1~��C��YU������W[�sD�Іa�\���I���l\�Ww�]��n�899�a	D�s�</[�j���
(��=@�l���=�[��U�^,����A;zd��1��B�U�"Ms�K�ȧ3mh�F���$>��oy/����@��]k��p�<�2�x5�B�gF�7���sk�1
�q/e{Cζ�Pm�fC,�Fc���Lx[����7s�����{g8��"D�"h�3��9U��i��6Ae����v��I0˱�ɢ��DE��� �ЋZ��7�C�gn\`�m��%��
���V���s�B�R{x
qA�\]0�_L#�|7����o7z,�舋"��S$���h%q #f�>�, ��ԇ�hRF�!s ���WKV'��>��b�lT";vX�#8�Ͷ�&������Lp�ٷ��c�(����4��1�ٳ��S�ڻ@k��GE� q���EM�4���+��zƍ)1d�$j9x���ך��`�ML�Y1�)�&\��Bo9��>���s�hy(��C.'˵�ֈ�ә�^�T5���tk�������w�a�(@ �＀`�Q�M��,�� b���ot5���/�$��������������a��J��سe���l��'���;?-�j�N�X!��Ъ�1�~��K��j��.�����	o�:��o�-t�����o��j�l����
����u�L��|�[����0�|ijtޮj.���S�T
���_�M`��-�Η%���M��ہ�GÍ�l�B��r^�7�s^��'d��^ה�`x�+?8HON{t	^t֎8j���s�)K6Zt|�����>�9���E���K�^:I��r�ץ�^��>��]�ټ�������x��Ziϥ�s��M��y��m��wNp��|ۦ���RET�-���.?^zq�㱎(t����.�<ր��Oʖ��ޗCWgM�6Ӛ�ji��<V�ҭ�Z��Z6��4F��W���`�w��'�'������7�'�������}������u�z���v��ϋ�?����u��>g���_������>�s�y���}�_�\n����(vqPc��PLt�g�}�b9XU�B��r�|�=G��>O�x��s�ws�m�x�+���#��q�~�Ρ�G���b=/}��э�_o�<X�����������|��4& �T�B��;���|���f�����xRכ�>�p~N�Q֡`�'�Ŋu`j��O���ۮv�*�ƴS��$u �9患+�����;�,�iĤ__��S.�����[o�%��np;����,Q�Ƅ��w��s >�AjN;e#�^1�SGN��/	*��Gj�1��2[cQ�"m��<S�.NQƧ[�.F*���\�[��U̟�@Z�&�8���bV��8t^�x]q���S�񏻼��͕�y�0I�"B�	ƨ(o�?[��FjF���d3�n��9��Hi�T���\�D��\d{#q���-̸�z�TK�:\"��oa�Q�{�k �3��m+��?�榒f:���wH��%t��q��fL�d剼f�Azn���?X�[zqn�i�����d��z��(H�ʍ�y�\Vߊ#o�RNn۶1^�:	&�.��4�n�h*��V<���v�h^ĵZ�sy�;
*J�K��k]9� ���u�vֆ��\��B�%�$�ȡW'��Y�ȝ�F��1��
(�!w6p�Y��Ǡ�����I]�Jb���N�� O�����ʾ78�-��B�{�~ˏ��H��e���6�J��Dv�V�Ff_�ZH�'*�l�P줧�+x�d��bJj�(���s]�^��?�8��7���J�A}��&�2$�8�ݷ��?r�&��EUZ��
�t��6��Ub��p��uܽ��leHJ��a껹��^�zYP���ղ�7˥Prat#xU��.���6�V���]��F��Km�I��wG�����T�N�"zv�y&�3�H����������DQ ��l 2�}�T�Wxl4�L�q�$�^.py�2����F\��UFҏ(a5����1��OE�<#к���i4��H�:`@J�1oRw�3�PTd܊���°Ӂ7�Ȏ��%�Kz��J��v�F<S��c��]����1�Iч�ZP��B��67ņ����8Z'C��fHN���uV�f�<��l(��.`Glhkϱ�P;���c���ρ[zd��:j�e�=I�K����5tL6��{ߖ��W�w��������vr�c\r�\�js�ަm0���$^QD#(wm�s��M>y�XF9����+�m��f���^Aq�N�_�+��,n�{K�0nR���ei�8�?�L3e�)$V�x�Jb����UIe�nm%�l*NѺ��MK��w7��!�}t#�����V�xѲ>�cAȤ��l�:�׉�D̼eCJ�b�B�m��.j*��X�9g	�N�z��׶���M�A�;u�eX�n9�D�=ï����<ċ�djo��oi%�R�D� ONӌ��wM�,�8�u~Fg9�I�N�V��j�]Y�: L�n�׵�5K�k�>����4\�38K����`�t�aHɲ^�AN�C��h���ѵ�mU���B�[t.���,ީn����
T��d\	'D�^�\��M+Az�.7�s{��:=\9u�r鞔���]��qKjzzJ*�K������aU?�=�;��_G�����?�W�������S����I�n����F������:l�5۷������KM� *n�j�ܪ:9������6�x�p���\��q��I�!�UB��}*�:�a�fw���w��[�
�Y��sp�i�Ģ�s�w�´���1��G����s]w@���u��'l��o�Sh;~-� ���O�>(��,i���|5�����U��`�q���|igp&3�̦�ʺE�~�o�jFr>X�LT�v�+�V�ҍ����x�rˋ����Yg���JG�|�@Y�@ 0�p��d��tQC�w��u}�-5"�o����y�P4�q�����~��r�w��w_��ws�{W���^���/#޺��<��>'y��K�v���{�+���^�����}���=/���N�����I��c��_��<�Y�A��-��C*�*��*�����~]�C��{?q�n���{q�w={3�Jp�k��;�KeLL9��^��	9��@Q%������|e�ګcb��Rv���?B���@q��������M�5���I�4~y�j�H�%�2��9�2Na}?��I}�5j��)}Bsu�?k+i��NZ4*�bM�bH�u#?<�9Ԡl��Qn�t������D����]1jZ�{�{f3mc�Y2u�9f�k�H�ѐ�*��v��ʏ-�Y�񐅳V�<��l�#�Ep�;#?}�$N7%���]Q-��B�@�HR���o������Y�>���1��?_=�������{?��\���~G�o�7x������_����}_����}/��_��������t ��p %�&����خ~@4P˷j�c��.`��
B",�$�����)��O�sG��%�#�Y� ��A����i:�дC��U�7�T�JZWt�(����uG�������ql�Y�@��Ts����cl.�f��RՕ��Y�,���������K�|��@�7�|�M��Ҹ�>N�����wo��G�Q���V�˭f%�I����6�5�:�1� ?�`@0C��c$����A2T�;���b+N(�1��x��� �
�1*����>������y���q��ױ�u��c�>/5���~��~O��_��~������|��z_��_�$�9������-S������{��� ` �t�X�dU	�����\l�Zg�Z�������"�Ѐ%��ֵ����i�T����\gB�̄.����w��9��v���yP��7哎)A}���@�wP6�q<PG5����	��뻉�"��GB3��#����y��X��7�y�X��F�G"DZD�od1*-4o�H]��;��ϓ�ӀT����?�+���ڍ��}���c��'�Q������5y��N1~���N?�>�S�=������_k�l��n���{��3�:ё���;L��C:I2O�
~�<'�7��!�7۲����/���5�P:_a����g����w���%���Cǧk�On�2LϾ�3 ;'�w�yP:�N�H-��f|���Xσ���K��-A" �dU��$Z~
�h}��{ݏp���t��\"��_ ��o�?���D�e�l��Q�b�ao�j�
="�	�����M��S9�tj��&�����Wu]��*l�6�Dr��sDDPD=A���r��m�>��^��%+���v��V
')&�~Q���/�?OP�A���x?Mϥ]���3!6�?�AQ<���ڮt���
�u	R�9�k�#r+4��3ml
������5����kh�j=��>IhZ@�X�?b���w� �/=>)%|vp�t�,�y��������d�r��IU��T/+���H<�c�7fa�3�H�T�4^�}�S_�Yă�r�'Ǟj��:?G�?��؂S�{G��w�:zB1�}0>�p�}��:L�xE�5-�ȣ�y�=���5����������0y��d��-���Z	r��F���m�kDG!J��"�$:���Ld��'<Vn|�$�i�me`�5�����H!�@P�b��w*���QMMn��E��̅�Noa'���vᨉ���w1�ix���(�\Z���ѥ�؈Y�0���mU:+�� ����1��QN]{��44���P�.4)?��{�����=��/X��~WQ4��@��&L���#�~���y�﮾#�� I�4�"=R�����l?���f|�j��'J31�D%Ԅ�D��������"E�o�@��v�<�ٷW�n�{�W��03<��^>e�n�>`����B\Zh�Z�19�����X�>�p{�-�µ��ߏ�ƣKs�����~1DzA�P������P��)44�Sn��{��u��I�{B�r�|��;��W��CA&�5��W��`���6�?�հ�͌�g3͌�|��հA�S�U��5%ɬ�Zݔ������!I����E�!\�g8�X�Vp������IfvNokd�|Z��l�`4���Y�3lݢ�������<mʴ�aUT��:;)$h�E�)0�[��"n���:���C�,�b�p�P�R����X¹ڔv�Ԣ���mw��٣�n/�."�#�4k��F���	 �<�3�Q���%1��h<%#
F��+k���#,�fA��{J��j	��Q��I���p�"�!D�L�5F�w�U�WU䰕pce���E�4
(�y%���ݷ�/bt�-��&'Z89�SV��i��
(�s�.�Ֆ�5�9�XH���{c��i~����XV抍�ksu�`�B��b�&X��b��J�� H$�����p�Щdkl�|9y���	����sYxVByt�S:�Ѯ�-�&��{�����8E%���}g�����j�l>��3��hQ�{��M~Mv��j�ԣbbsM?1��E�����ݏx�O{�L���9��������f%�!2�ۢ�/ii����=�C9ѕ��m:�]~�Hߒ����&8�=��?�5��B
��]�>��y6��$��q��jv��T��s�C�'��j��K '5nu��!h�6�3��8��{]�����s��.-[��*K#�ϻ����LJ\�I��8�!�u:�8�fY#�o�ѝ�ɒ�EBΏsru��Ҍh��2���d"���1�$jI�/w�LL�n�2j��͍��I�M(jL�3Q��z�������1\d��Ux�c)�1W$1��8�Z �����φ9u�E���E.un�6u1�| �V�t�8���7�ʫ:��V%���T���S/�]�]rFTg��q�i� �")w"�ir����pB0ʢ�����?�����i��LѪ��y��5FA0LL��ɬ�;FF��K���m{HOsT�9��&���V4��(��@"KC��c:�E0�M-C��\�$�Q�1C�%3!�ud�:��td&�@j�S ���$(��@�xy��k�3̜$W$(_�ݖ�lw�E���$ʚ������Q��19��w]���l���3����"�θ���Zœ�"������⢠����b.��Tc�mW.����T9ɡ�4�L`s�.�S��%(*H�V�������c���6v`A��RRn��q9]�+�;�jj,��1R+}�s���rkƗ�=t��	�L���9���:rt�2%Ȇ��F��Q�J�G��H%�+JX���������<�sw�4������$�#��K�6Z
:�� ͢�1X�l�1@�>H��9]p{oeq����.w�:Q� �G���*�a�|E�bn���o�*%�U�����M��� M6��Up�#���ق���R���Y �=����	�BLMj���i��� �}G���_��4���	H����b-|��󵥊A�@Ȳ���u����p)���#	��J��x2G�$�8(�Ƴn�&�坐"%rt�a�Z�#;�1�����
�W�g���*�V��=�lҭ]�l� d�$��N�\�@��s��a��$ܲ�� ��\�5#��V�b��i䙮��ZL"V �crH�陈�$���fh͈�L�܈�$�-�Eٷ"�\����h�¢�P���iX1v�0 w�*�Q6HK�jC!�2H��� �]Wo�XUΓ\H3{Av����G��S�%��t�o i��D��:e#˶�L�j��Q��_�8<�!�B"K�RK"N֏��Ӹt�0 �!��n���G9����a�Cq�q%��#��S4.�3)=�������a����u[�T�m�9'�z�jF����s9�8pd2,$N"M,@H�PPm�i��Q�z!�B�:qFa�;�ZҮ��uZ�IB߿SF�ŗHpk�gteT{�Y �j��>7A���8���o�U�Y��!�G�_���`i�Mzw�P��v�~m�(����-�dN�PDJ]��;�o�A+*��)2�Wѽj�,��T-(	'64gRH�6r�?�"��ǃ�N\��,J��Jք��=o��!D�Enc�V�.���_������&&j֊���"��"\��r��� b�BIܹ�آU]�b���l��AB�e|�b&H���:�6�(�Y��d�If�H��,�nʻP�RA�Ș�!Ctf��R�� /|�^Q�(�ؒJ�!~b���#��{�P�Hz���e�2���&؊�iҶ$ڛLX�3Z YT�(��Rԋ��Z�h�/�(�DB	%�#6J*��Pp%,�b��Ң��|��"lYJ-�i7,(���ѡ��fFIj���s�#�
T��sL�j�VC �3aИ��s��D����)�I���<a�0Zmj$�Թ�G\,������$�&�/>~~A�8
$��z'RH�������Ȧ0K�V�6����tL�`IW��R�"����H	g�al2N�W���|e��aK�3(�JK�0̧�zF5#r	��E'Q�{���$�a��A��d��u5@�L8�J�hLPN��Y�o�ںB�-� ���'ߐ7�8u;���'�t�����p�@H�&h���PBLUG�,h�$��9�Eb�+7a�C\�b$�ڃ{� �����0f0zS} -塬$I)�.d�w(L�̒\�B	%��r̎&ɒ�f�&@i�&�lH�X���0O�MB�xH��G�/"Fƍ�Q�0�R�${�G<�
 &�aP���^y��"�rET�%�,B`�{�Er�*�0�	(���w�I��Ȳ¾���T�VA��������C��4��'��� ��5H"ȷ�r.
fqB�@J@�A���僞Q�cR�0�ɑ�թQ�l�kEDbN��!�h�$7�!�(IzT8�o
s_��}��+�A[�������F�G��/Y 5" Ո�D�
�>���$H ���H���-(Ag�!�}^���)�UB�ԋN�k���ُ�CH��#4^�pWY�iG���=t�]Dj��Vj�xu6#����h͚�Y�s67�b!B(h�,�Hkp����$��7��^$�R���:y���&E�d!S �Α�賑��L��(��	=���(�J���d%6���F��-R�AT8A��	������yA�*�-��F�����fA	2~hApg� �túd��1�8ADxz�"tj��9���^3��n�h�c!`r �*�IAw�����]km �$@D�	�38"@)�I�(�
Z`�_앧�)HƐȺh�j��t��8@�93hEcV�Z�'��;��H����`�_���ş�����ʏYA�m����e#Nף��nRh�C%S�����.�I$�H�D�YM�z[ѐ,����PR!���&e1�.L ��DnEh����D���Q�RQil�ǉ����I��"S].��)�ށ���%+���d������Cl�:T<�Zl��U,Y��D�&�h�B�P$�[��9���0����$�`�~���\|~i��0Cvܨ�9bേ�ڂ�К]B��#�k�N��p9d�@��H�ˢ`����]�fZj�{X
���8�?)��:�e��$]�r�!�
Ũ@$"}W�B|�����?)�Xτ���H�Ն+4U�[$�H&&B���֨��5 �B�ɢr��E��0����I"fkN���B2{F{��T�ZZm���ܥKȺYW�eJ\��j��($N.1BZ�.,į�؄!?�����~7�p�x�ZYk�ײ�~><�}�����DN�rl�J8��yhFT$4">�c?��ʎUF*���^��^��m���('4U 8�FIV*<��5����=�&a�O�4����}�����"Ъ�]�����&��)�Y�N���Vm@A1 �ť�&�[:0g?	��z��=��|s���O�P�a$��)E��U�Z�bLQ��)2D%���]P[���И+�B���Ӡ��H�hKAQ#E��Q��:"	 ����$��h�$A,�
�TD�cJ9(����bR�f�}����F�_ �S�&#C�L�t���viX�폟���HH�Ć�g���'����:��@���~��5�A#��kǞ����&I��6?����������0��0�A �����K�Tk�
� �a�^�SO��!$�)E
ǣr��;I��qɉ��$2�#V�:E��eF�9Z��S	��/t�h�D����"�#��>�F/򼵚�W����h]O��R�h!j����,62KD���2lg�%}0�C�S���R����o���:8LX�,A2�PdUZ�ڬނ��)U�H�
GX#��\-����m2�P�($�V�Z�iBQ�6���<qt���Eh!�G���۾H�3����FwKS�8����iɩ6�桸��~��[V((��I:�6tβ6�؟AAu��S��X�bwTDfC�6VT�m�߱���{�0i�R�Cډȍk�.f�l��6�0#R�d��Ъ �QVN��a9�Q���{i��2Rd��Z*�J�j0A���u��	��{[��I���$���G�I����e����$$C��t�/4��C���{�}.�h�'͢���j�m�t�F��4g�j����&#���b�+x~.?���*���U�\j?T�:�1�7iЫ�Hb��] �R~<��	j���4 ��!;>nG���OF4����%����QzBh�DA�e���ce ���fB�|=�'�۹�{�1�Я�z~ğn���h�>�0��`�$kR#5�W �ȅ-�,�J̩K��ԝQ���\����PJ�(��Z�mP+ʙ������3πK��4zJ�X����q��^}�˭2׬ V���R�qZn�
��1x5ao$�E��9����X�@V��8ߪ>���C2�ci��g���/�̤�i{!����J�L=�#:�"C����� �
�O��q~GȎ��U9Ɓwk����:�)��V��kPNl��v01qG^�F�s��*r[��B��b�8��I��~��pRü�l�J������Ȉ�ٳd���^��;vZ��>DMi�߱�šs���SR�*��ȃ+���R��h�7p�!����[�*�&*�I����3�ύTZ�QY$($�yB��Z%,ԭ 還^Q�|#K94k�Q����g|��U����� ���R�(%���7����e���Q�M�k&E����j���U�Z�Q\g5�j�T+�^QT�<Lo�
6��ݠ�U��S?�������%����l�L�n��M��9Ԑ�Th��R��Ü�r��T�rV{�����\�}G�D����|)����:�%P ��~ʶ���@�0���iR�I�M����Ťh�oZ= �W�1�q��H�����/:*R�g�|iJ�Pn����|���Y���A�jUCRj
� �\��bR���_��}<T{�SWc��[���-s�r��6��-b�:d�թSd첊�a
J����E�U�rE�H0�>�{��F�M(�M��ISI�dhxoIH�֯�9�\�<,ؓ�|?ӵ��"r74G.�����p�+WN&��j�h����%G�~����������hw�Uv>��30{�d_G�޾s����`|sJFUVsB����M��=1����K��0�+���D�5Z���������<l�M��4�r�>���Da0�g̉��{�h�s#\3�+D�id��9N�Tr�c!5<M���s)gT��f��ǟN�t�m�'HbWȸ �hlFRh�oߥ�ϻ�bX�@�����C�(fp�����;��^��?C��R`������ڝ����3���"�}�sPr��u��\L��&|
f傥C�ݍ-[	D�!fXZ�ʗ�Vg+:��zR�ĊU�E���f{#[i�6���so*�!!J�ŧ]�殥�Q�ջ�T�ڹ����A$CHY�{^�P�9E!s+�%�R4F�a�'I�Ѩ���CK�]�Օ�|�;���%�k�*�q"�Z��'š�$.�4����YT�JO�{��KE����yT�4���w�$ѽf$D�B�@���[�K�$���\5i��mć'�g:2�G-���P"�^�K�]YFjWj�`�tU�����~N��%Pn�llUr�UG^��G.9�DL�Z���3%ֱڙ��HV�������[+X�������+��KI(����y�YewRʤ�T�� �Y��S�t��d/��5�E��{R=�
��ckb�r�Uh}g9!A9�"*.�b@I�U�pI�1d�CBW8���>�ֶ`���e���H� M��MZ,�St��3�7nQ�"N��R	�X�\&�
e6���nz��5 �Y^BN����pJ�mI9�A�^�l��Tɡ�r]�X�s���C@��(�f�?�Y�R5kt:[F>�
r�<� ϭ+7���4&|��x��ak�D�dX5	e�	 ,A@l��L.���'W�B��
U&�Rn{�[��[<�j�V�r��Pu�cmVM��PF�Q�����,�a<*���U�̿0fA��[�)�N�q",&�Hd���&ٳW-C�QL�J��=�X6,A4I�D�x�B�A=*���EUe(iQ>��k:�m�L,��J,-�<:��/I�����b�I*�z)=�ﱵ�X�L��*��J����e<��^������U.�]�[��7���m�	����3���C#��Tc��@��qA�J�#��Ca9��N����"A�/E�H�)�����$D�7 k����Xۊ̋8ܕ���(����oh����B�Q!%�fYHo�؂��V�8���Ό����e��6 �;4��hL�h�#`�T�A���%�U�"M�RAe�)��к�4M�V��Lp�jY��έ����EQ	�hj%<�1ױ�`P!Rx{FC�9�9�5tڴx�R������+��'�N���	OG�����MG�0(f�lr ZxU���Ƙ�f2�7*�A)�u�����faU$7�~iAV'�YZ\T�ef���2vkYXՎ��MU�!ş>����}1��Ld(�7,����!$�K� �r܆��SI	��;��4�rP Uj���+��S����I,�]|9Z�j�w���"2�1�p$ͭP[rlBۑ���f�$a
	Դ���r�'Y�*	&Y��b����5���H��P�I5����&K�D�i�4�6i| $f�{�CCAdvR�� ̦�;$i������r�aE�*}p�!� ���F!V@�c�&(ɝ��N�Ѱ�)|�g �nO�>�?9�>>��$��E�i��3Ix�d.'h���L�%9�������{�4�C�48�����U��c Y�I�a2�[5�4JA�L�.�nMڅ��_7d1��(��ׯg�鼩C̋�D�n�!���
��Y��1d��ekZ�d�ɰM�Z5�:�ZMfK%l	Ѕ@[Vrs�βI؄�8�7��ˌҶV @L�,�2B�1%�B�2��UV��_]Fέ����&�(�!��K,BR,"h(����Aʈ]T�&�Ej �L{D���4�^6/�����7�^�v�U	�X\��Y΄�2]o<����MP
�Z��ߓ�HgX�mb*�Il�&4%)&���]^	s�cybh��z�U$�$m ���E¤��Ci���4(5(�5�t5����q$F^%�s��`��"�C���.֝s�H� q����!I$Q�D8ץ�1A!q*
qmE�~'���PFF�l�(ȃ���:��zA��a6���U3jbU�5���B�by�����v^'���A#���&����FT� ��1s�mT��R$�A�e3屆�y�B����"�X�#�A6S"
�q6��"��E	�e�4a$�	%���Ӕ&#:0�� ̕����O��_��!�������ˈ~�='��4,cLK\s�>|u�K"X��5/@]+BP�.�'b*4�P�
VHX��˿B�IMn�6. �I������b$	�J1MP ,�!$4��V�Xl(����̲��m&�+
	V�{\H ��6�;����Sa��a,z�U�l'�Y�[Z�d#�6�hi�����z�1&�����LTF$H	��̅+)�L���(�5*[Z5<]*�%�3;�P�H#(�@إ� @2!7�(]-�Ԙ����C�5kE�J!�$� Ü�g�N���l��Rn���򾱝(�>��D4!�|J�c�B@��7��44�H��q�J�F١+D �IH�����¢�I�@��f�ՏM3m���Z����!�5�o��!#4Y��TQ�p�s���9B.ە���^�@��E���6!�)���,��MA@��8�Oe��i+�Vt-$����Ri���e���j�B! �*o6Zt�BD�$�Pࠨ��Y�].ȂrL��Z�R��T�W��@�Eb�ؐXH �%0os��`��������7Y�E��ń �d�#��D�#D�!T ���h�,8� ���`A%n�v�3'0< 0&�v�V�(�Ae�,�7GH�>"L$��%k%HJ��P!&4F�eA~a-5�����4b�`B�e5JN�h��iړ��n��5t0���*�kjY:笝0���V!T@L�L �`Q��F�L��T�U(�#u}Y��^dd��� �� �PL~���C��T1�I
j�._y𱦐d[�j>ۣ��B�cc�@a��>��H �|Tg���������!ԕ�G�e��	m�Ƣ��d9LR�D@��H�m^A$[Ec�R��T�R�Mj�c?����_J�I	~�L��>2$�
��:�4H�_{�D�
@ai^@��Y��{��4@���'N�H�TTrU\�s��Κk�]�
��.�T�P�_�m��f��KY,�]k���Ɋ!�x.4�h�R�Y�<�]�<I"~�D`?AR�_j0~_ھ׃ �"�T�QeBӄ�;�h�P�B ������ЋQ`J�,D�m��I3Zd�Hh�v�I|��et"�E
�Ħ�(ZA���K*q���4B�Bd"�j��,�&O6"-�U�-�i9��/��b�l���RODJYNF@����\��12/�|H���i���Ս��~��&h�Rj��)���GX�ڍ,�"��]�S0 ����\�*ǉn�bp�Tt�A�D(h�{qY܀,$�4b�Ы�y���h�2��&��m+8ZvR��¾Z�hP��D�4�a�A�B�j?�k)f�)#2�)��f�FD� �؉\��$R�$
0��	��"lU�/z��8���4�z� �-T�f��/lM ��F��
dCHN�tC���D�T�"E�f��T��!$G�$�LҰu�����#(���,�`_)���Z8�|�8{��,�1aX��tm|�ȖV��3�!K�Q��!�r�}LHk�"bB�(%H���@Q�����J!�Q�
�i�Q��+�L�����eG~tq/!_d���{�?�,�@��/��v���J?K�{�8���H"��3�_�~w��-���)�=��v��|�������H���v;�J�
�Ԃ�3�K�he/�-Xh�DB�Ŧ%�)	A�B�{�y$�aP�)J��%|DZ��	a*_PGhB�o�Q(DV�B�:<8�PP)G��r��<�&������{HԐ�#6�E��yǿ@�����	�"[��ϟ��3o|��V�Z��3�񔍈ie�9�A���[*_���9��1�Ii�\P��j5Wڑ�$\�V�$0�P��|�|��"��#�����o>w��U�G>�������4���HwW���XZEU�$�:	�Cd|~)���
-i���2���Z���J�B��O��SOH����7mI���I:XH�#��W(F=HBQ��!ya{ӗ�7��,��)�E(۸ټ��,H�
M�Q�K���;��$E�����L�&BФ��aj��li0�)����s .��FG�o ~�!�w�M�壜� ��9))(���������ڧ���/��,(�+HoJ������ �&��r��S�ԒnM8������T��1մ��{���KJ�;7��&Hq+P�U��'Ϗ�=��z��?Ŗx��7�<�����p��޹����+J�~3�o�X�KHh8(X3<�;BQ'X0��p��ݾZl�t�����9�֍/�u�#eg���Y˙AZ��<5����=�?�
��K�28�xHQ�z�~ע�t�8`��������ػ��M@SP"�� B$*
� �K"����
0�B
�m�~���˜�l�Hn��0����"�(�H�������~�� e�MB�`%w�h�IBaihK?3�w��������lP���&��� �dBQ%IT�BU�%B���J�i��
�
�( �|8���MJ��J�3�^�h�]������3o��<JCk�@=����sGg��C���en+�_S�y��=5�v�8
$m��I�} �<���tځS6P��F$�
)�=���b&㢸B@���$0�Uo�Or���ա72B$;���������>;��T�Q�
�\�N��a� P�$R� �}����?`�!�u����0D,�H
��{�K�ݗ��@������q�>U}^ۡ�(VD��7��ފ
�.�}Wo��z*H҂/��"�xfb &�64T�j�,D����Y ( �>(�̃�!hڀ�`( 6��໗p󽧿m.�'L P�a@�$z�~�����G��;w�jQ75a�6����	�{�H�������ݗ��Mhp��Ez�8�����"@��?`�I�~��v8W�>^i?�� 5L�/U:����Y~I�[i~�& (B4 B���/��;�Ws:�x��v���y���7�yO��B�ҿq?T=8���=O������.&2>w=�s!�f�Tꀐ�{'����k�>���~k����y� ���n����?��/���?��~������#����^	˙~��N��f��؏!ս�j�ܾG��]�-�Pڐ�%I�z�����ܘW������
9��r='��WA������oz�����?��^R����a�$&���?)���=��T�9 ��g��O��\?=���z�GZ�9�)����8��~G|��"}��������=7x����:�{�~BB�A���N��u���}����}����L�
�(��������SX�U����A�
'��n�_��?Rn�+�Sڟ�V]���0��v)���?��w����
 )�|�4Mt)�N��(���}���+pt �\#�y��s���e���+������o2zt3�j�����N��;�cS����{���J:��0��m����"�����ϳ~$u���vz���4"<�$�OrO�z�G��������_n���'���|c�d����=���� kl���Ok�K�r�'���f�k����JZ)��p�@4���� y�u D�KS$��O5����cE��Z?��Q�ݘ�nc���+��0W$�eZ-�%��S�3\7wn��\�e��Q��&��B#EEc�(رQ�4m���Q�4j�B�5&�Y��#D���~[�￹���J����wE��-0qI����#H7zxQz]8���I�14�<!����3��BI�I�������w��ן���o4h��Ad�F2v�?%Ttz��3O�������O�d���a.i���h���K�9�$�"N������!�mEɦ�u��f�"�n��t�wp���X�	�:��~���&fI7�c$�7rK�1!BP�+f�f��ٛ�6{�Lƹ$�Zȑ����+��:�ֹ�O�����d)��K2+$�d��3̵u���S�0]���JRwk�%��4ddI���up�Ū�l�IL�R�	��:k,���VADT�L��n����sS�ݮ�wu�1��NwN�v�]��2\��˝�wuɐ��s{ֵm�{{c^����#�ݒ�5]ñr���z�#yܕ$ �		Y�F1qFK��u��u;1]ݩ�WLc	�̐�9������\74��v#b1�J���	r��Ac1��(�@�	�#���*�/��G_�W�j�����o�:㻓��~������*���8��X��;Cv%�8+���)��"�ᶄ� � �D�RwSv�VEF$���
8J
M3ek��$)mJ�� �)@�(҅%����BQUIjJ�+��U4IdS"�XC5BB�5Qʬ�-�[�;t2�T�!X�6��T��X�d�ȱI�d̙�d�d�������u+x��J�iJe%c�'��!�$#(�$�%B�1T��[6��"���"""��V��TOf�w.��n<۶���ז�`�'�S�vg�M�
��j�`�b�⤹w9��������d#A�ɺr]s��t���+�k��^�\\<��������Y�F.�0��	��#Mt�%$GZ�%%� a/������{��Be)))����"l�$E¾��O���x��[���$�,��!�V:��3L�C�\�
X�m�Eg�L
G���3������p>�Q/� b�&�lnI��\	��'�~H��'��N��������L��6O\�_�;�;:O% O9��9���D���!=拏$�SI�Wfq�ɑf#��eC��gb_��|@B��cp���*L�8�7H��ݝY���@�ٷ��;F�hƆ������nT�"(]ݙ d[�ܝ{�Z��Y��$�wdpZczuC��E��$��a�4��"�>YK-�7��&���c�
 	���D��3:|�C��;s7pP����)ĒN���&y鄳��.ZnjW2	�8v�p�̜�&�K�F�Kp)4��.B�>��lՌe����5�j7kX�4m�i!��g�F�4��5�N����Jsݜ;pnF��`1���݇:�٫o4�2ƺ�@@̄����ޛa�Y�O9%�HzD�'���c)�>}��;$��	�Ԙ��> -�dy> L�r횗 ��5X��v�2�o-Fc��],�9���ϩ1�d�w�ܛ��KIs�f�$۝��ld�I��F�>�͒�p��HDQ��x��!�6!#'9>���%�>���л�s!!���f��ϓf�$��k��s�ȿd,�d>y�&�,�7#��̶Xف	p�]��������sr����0��)����I�<Y	L��Ɛޞ�	�	>�=�����d�FHv�Yz�d�����f�y�	��@�$ʶ)������(�+_�����$��8�5�0���@;t�z�����8�d	v�lsƓWL�i9Ԇz���M�	���p��X�I$�E���>x.~��I" _K������Q&���rJ7mv ٍ�$�.��ح�M�t�o�N�M;2�XM�L�M�j�he�$�f�4�Ba$%2Nߣd�߾�}V��܏�$�;(r��s\��,X
�Km����bD	-r�,�o�@a�����#n#<���Ðɹ�e��5��I��d )�`�ßL��7�م��y�q�8I��}���Z�K�ҹ��2���6XB,$A�3��|II%ȳ		�x�u�-���B{�z�d󧝓�e�۟	���:�d�trd�@5��f"��* Y���4EPs�Eq��� �����8F`0J��g�8JR%�Ep.��^ ��i�S��8k���7M�j��moݭu��(�y�UAD=���N�ӔmX�
�n\�wc��Eӧ]�pRuٷ�!��y��W��ѹr���s���[�r�F�5�mͮ�ඒ�i�v���oSfLĤ`��%�=
LPoU~?�E�ԯ���-{W��"hF�짮��t8�FP��
hZr�ōĮj;�lTUW2J�"jdS�0�a0�d�& �He\a0�$0� ��`NGh�ʊ��x �`�a�{~���A����!��o�zc�����7�"�+F� �9�k\�Ũ���lV�mk_�mU_D�wE�4��3O�	30:�=��=��o�|��ϟ��b�F�RY��#6B1�"��EA�wI����`�U9��f�a=���~~�4C��J�J#�����Ҙp���;=��4 ��������R dGrP@Ziuu03��d��q?�C�0l@�~�Hp�U�S����$���J2rO���ɘ��z���w1�����>�`���1�\�9ߤyz��x�p/rI�;Bd lXA�� ���>A'��>ß%�|OC���A��=a��#��I��T��<g��ft�հ�����?O�j]���c�|y����'c��?�W� ���t��h3�X�*�GɅ��c����r^�Kj1���ɋj�/+vVצ��)���0�Dš�y��zY�J �b__ԯN����I�d������y x!T"A
Dunce��bù��,M��'�f��'��~��Y���ݟR2	"?����!��+	��� I$g.��q��-22�Ȋ�m���PC�?��P��s��	.�F!
>"|IJ A�[~A�L%��d� N��2@e%���=>90�^���� �{Ns](��4\���9���U��:ȆU T�	�y�}svi����	���2��*2)9(6X�w_-��'��U����})� ���8��"$$M%�DX1�~���{���R�����  w�e��k��Y�ߢ�h .y�k�$:��n(9��'�v��y��2�ǥ��i>�_����w��;^�u��a_|>���F|��z���Z�w%ZPR��Y������ܱ���v�����t��*Gi��d�_Yz������M��;��K�S���?{�x���6�R�pTq�Ο𜛟q	6tW�wlZ&�_�H���'R��8FBw�a�Q��X�����sh��w�{��"�N�C�G�T3;���;�T��I?�*��������텰�QQ��Jp��P(biy�YQC��?+�>;a������	����~[�ܭ5p* G������
�9�lꉾ��ROt������ �_�)�~���߃Y�	~o��w�����.�{�3��K��.���ΰ�R��*���Ȣ���`E;8�1���c��?�=�N�/ ��/���O�a��-�6�;1�
��?� �=�n���!\�z�NX9�������P =;]x���]�B=�
���p(��@�+�_.�9��`��}�y������`bW����r�m޿�������~���� �k�G/��"j���Hv#������TtFO�u�0v������_��=v����������q|����~�~*��+H�D��%=j�0W�;wd�S��{��>C�_/����L����������G���ϗ���7ߵď�����O��O�^�4�?3����ג���	�D���b��`�������,�_��L~<G�֊<Q�^�v��וٹ�U�B���i���؃ҫJ�u�o��;�l�hRJ����~L�e���<���_���~�f�I��B�s�(��IވAu���o��G�Q�jv����ƙs�o�x�W����3`}T딝�p��y�2:А�ݪ�:�ᑁ�#T�0F�"ؒƊ�ZX A�(��4��k��P2�@}u � ��S�ʱM	2��`K<rM$HB^9J/'�sI���GCH�G.���#��~�+�Q%Q��L��H��p�����6E3IO�#�L��w�B6�jV�y�Dl�6H`.������vх3T�
8sI�@4Q����1	!�4m%)j����m[հ�f ��ʠ��u:��A�F	�אf���^�'�>�������"�}��9RWwf��ma{�D޽��q��t�c������A�|րCH���$�\�ɝ%�:̑0�e��@��ӘQQC��.�K���	��{eaܑ>��%P�Uik�$'W�#~��;�[���Y�Z�B��,��YFU�t�G`9��^0����A�jĔTA�GTS�N<E�s������r�����q�(����9�`1Sf��4.�0�$D��W4��B.ᶪ>�7υQ���Zj]�A�7�,lI��F)6����o�iA�'R"��˒NW�"	�P��M5Th�����$����{g�����&#�D��p�)%���n\�܌��9�PD�]3�r�����0.��̄�\)̃����8E��l�f���dLU�&�����7�	?��'dP�	�lS�qȊsjk�`Q¢���	��0����\!�>����Mbdt'��٢�x���'E�DJE�)P������-�L����ԙ�*�h098@^I���{�,��ߗ�M�3�� ;Z����Ꙕ�{�bLN 879g:KVXLCF+�_c���PCD�"��� g��\�A�j��f;�c�{*�0���x�
�p���L��o�Z݌W���&���k����¨��ve��ӊ;J 8����8��!9��N��2����-J9�95H�q�Cu�`jw6� Q�ǰ�:*�����8�@W��v���/n0k�h�!)h��)M�8�yI��� �P��K�
Ȩs�)���^��'�f�g�����(���4`�o�.d�cʊ���2�|�0�6C���
��45p��{x�oo���}L��E(Q��%����U"�`���yx���4WB]������E�\�cDb1�\̆��΂E$�S���:��˺��sWg!�r]�]�np�t��:�b �5
%�]ع�rwvL��n��&l��jP��$��j�x`5��(dT�*�Vh�
$Ⴙ�m���GtsD3 PyݥPz�<��2"���R���~N����fb�N(�bʸ��AT�	���EQ�e��`Q�͵=��:S!�w�!j[�3]�M�m�yPv��������d˄���a�����0�:�].Y�d�Ec��o5E8]X9125�Bkq 1�t���h��mI��AL���c�'V<0�y�9��[��.�� [��/�]��
��XMj ���f��(��§&�`����GG���k12'�]�0{�� ��H��,�\7� ��01��|��`���o�x<%�S������+{Vb��+���QReL(�8�!�� �ei S1%�y����Z�aX(� X��J沶�W$M��# ��� ��	^1�\ 	�FCX����h�����8A�xq~#����<`z�8a �~:#� tW���T9�T=b���wP�ǀo�M`8z��G?���+�=�E@fm�u�����CG�9�����&^F)T� �D(U�B���:�鼏 !@P��J��@�0�&�S�jV;r�����Q4n�Ϩ��n�r�8��{G$c�3����L�B"&!٨�x�yǑD. ��y>w3Ft@�5�� \�PC�6�#��ڨ:�5*��h�2(�h�C"�6
���8E6r*���pkM@��"�9�Z�9o�©��J	�������<`�?o������9 8��G��2!!`	AFU	R F9U9`2���(����d�Q�M��@�GL��6��hj�OTz��=es��C鬠�#)�^��
�W�=>�˥���yۙF��἗����u��yl}o������s������}�������x���p1��y��L�"��P�nT�*$|�Lv�Y����d<Ҥ8��T���7 ��y8T�ܰ� t����.`&�B��
�J��.H�������`��OC���9N<2���S�"�=�G���o��<e6 f�b:�vtJh 됤hD�5��с�ܜi�d���x������?l�|�f',	�B��@�	�>�90'#�#����E�@��u�<WZ"�}���N)�0��Wl��@�ªw}����	�'�s��v���rx�2�j(��2�v��h8 9�u�x��r
�"p��������A�������UIt�t�9.{
��dX��A�O�C���!����`�X�&����jؙ<�I���o5�>���_��<_��>+��?������=O6o�������������O�@��(�������?�|ȏ���}�/�<ɾ���$F�Y]y}_��{�u���|� e��J1��0��'x���M����?����&0Cp����Z���;�>#л�4�B��z*F|!�A"�����!�5j@,2���>��W��p���<>W�z�{�<���'�@�����s,O���3��/�?�����zO�3�0�_��� �#�������P�"L*�q���ϫ����&S-���I���������.(Pe�q�J��	H��;d ��PSP��%@�3>j�J�!"�~�1�1r�* �T�����%o�DR���_�	��gc�~�/U�^o�Ƭ�y�_�Y���ce�+�"��[/�ŒxrG�|$�\��:݉���|�����=��zm�t���������]غ�� M����R�̔�c��򥅦t�4O������Z�.&�?�G!�=����f�o�jCdO�M� �'�?�,�Zc��{��1����A3�߶ �f�f���j�"�P������l��h�o;Dd��9<���`�AǄ=Ĕ����s�Do�_7�ø.����
�:^�)�I1�~�2P�[
�$���`
g �H�٨�?��Т���'�}M O��{J����3�
D�B���:t�xOf�N�����Sz9�t�?P3�'��e�x�ɿ������u�Ы�\�I���-W��_��z�4��U���<ׯ,�'uN��s�u[����_g��ow9�v�:�M��߾���;[�d�������7f�Y���rd4��U�7���Lw�zw���j5F,EMD P�R��C&Hf�S5D�O�0dv�����,�tA1���
z�'��Z��C&�7���֮�&�DcF�m�6��z�Q��$��	
�����o����zoU�x]�>���>�}����=��~�쌽���5���z�(*Q�d�8��|hz��� � h�X���y���ո�����ո���?g���.Ck�����{lp�%+��.���(
��kaJ*�xC�o����*�( ����6���>��z�{�}��ߣٶu;G��G�e�oo��?����(���bx~�鿋���#����1��߭��T���2�֑�_����_��~�����k�
r�r�x�1~1�`�A������R'�VP�yE�;+ �?�d�����tQ��:]�����$a��#@��C��;���G�s�Iu�j���%^��ŏ/��,/��}�܇M����3@߫���Ks�v'F�3G�k_�#������8�[��?�=�#�)�d8��x��A>Kv����Xec��	�$*e���wCb'�;�M�!�$�E������'��7��9y
�r��3�y�!K/��~��>-�<�%�������v�X������z����}��~�%�4���p�_fâ�>���"0��̑,��Њ�B|��u��) ��L'$	_�!� �2Z)� (�`y��!���a�hDiEi_c��}~fg�mB�I�X"����A�Z��O��� �b����G���H Ц ���)h#�)kj*�������H#S�����E5{Ϗ��aS���H��wt�� ���Cd$B@I�}�����dx��d fH�@!B�*%"�<��/~��7��;��^s������}����O,C��R}/� �@���o�q�@�k�Ha�)2�w�����<?S�E���G�����?���~gݛ�@C�c�������C�_�+��T����I?�r�R�9@�O��ԠAD���w���*����'�|_���$���!p��ϥW���}��zS�/��?��~���`�~�����0�`��������A|���������"߈���O�=�L!B7�����ۢ~p���{�L�(������ھ�������<���Qt���9�e����|��?����)�D=�v#ƥ�ߡ����_��?��5|W�W����X�M�����}�`3�$?��_f�����'�6>(���ւd�b\��q�����W�D-�݌�*G@�OTIĹBc��[����]�S)	p��)��S�M ��mc�-%		�Tqe(��%x�Uq̆c!�)�"&^e�D���I@Z��dUW���X�EWjx%� DA�t���Ô<��z,H�S'W�	�E�a1��d��UBX�TN ���` �v��9�c��Y�QJ/�P�����)��o�����^8��)���8���FR�0�R �(PN_<�xɘ���������:�0��I�癩�b��;�~1�3R2������^?�t�������z���g�������ߓ��{՟��������~˭�����7��w_���P�������_/�|������p�?���n��?k����e��?�������������0*>��xo��[��]{�{��z�?��m�4�n���w�n�_���k�~�_w��������Ǆ�A�'�;)��Y��^��D�4�NE~Q�ف !��� ?ʟ���,�	�>G�~.K�f��@��oN��Y��!���'5��La�2>�c�uHv�%}X_! 2'�$�b�PV�B$�0�?���t ��^���c;�CV��_*������{��>��}�t?�|�`���O�n��;���{s�I/���_�}(��F{/�q��<��2�O�-3o�P�	��^�Zoy��{H)���B��	�?��+]�|H�b��C4��������kA��F��@���a�$3=g�K*�(��8�0u�R@W��m�R�	����e��CI��xB��~YH�4
����RR�U����4����H��<p�Ad�%k�LcIT���zOG���ǣ�Q�	_A�7ڄ��/�O��C Y�o���m݆�X.��X�mC��@�����?��z/��޻�Po��b}���o�!a�����R���7��G�_p�7���W��8~������ig<�����n^i~���N]�{b\�˷��C�\�-�n_������s���X������IEB����,e`Æ,c.s�Nx����f��w������{q�S z���}�!HW����,K��=�hA����uW1<@�������)L¤�9�9��4�iE�z��d��|?�+�|�)�d8:��?ˍ��OV��Ok�����!�	>m��2�S��p�����]	�	��+��JE��������NN��3l�o�xl��k�I!�w��~���g`IJt�o���-u@%�C�~ǟ�w���)��O��/� 4du�7�������T����#%C9Fe������s�ܙuRL)���,�fh�n?�d>A �;�ع�m4M%� I��O���h'�z����Zj/���A�D��Ә?ؐ�(��F	z���rDd�g���f!��XI�����#3@A�����ϳ���%�e��
E"=o�z��3=M�:R�Oȿ�44��z�x�֡@� zC��P�����T�$B�|��~ �5 }���;�*`!	R@�`$ID�e ^���h��|Y�H4�B,6��>���%�ӽf���d�h�q5�g}�.��2F^�ٚ%�����9q/�|c�2T!H�dYR@%IP�!XYD�����2����D��� ��~���ПsDs&�"UB����X�Or��]w��`  ���	��>����4T��@��	B&Q�$Y�aIYV� OH)�!)D*�hJG %����}o�;y>���L�2��{} �@� �R�H�U�un�����VqE8�TUb�����ZX���X�/ōí`��a�|� @L!B �b������[��[dC"K���r�=��'%a�!Q�3HPv�q��W����gJ�O3�^�����I�;�_��U�G΄[H���?�w����'���qTH�E�H���[ӫ~i��k���^�R���%RS`�ӛ��Z�G�����?����/�~n'�b�{
�j���l��	WL����i*3f�z{��.��[A�
�4E�Q�q��9�>W�24l���%����嵞�^�e��M,i���(�3���*��@�)(��
�2�J,+(�	@�$�B0�C , ���Ul}/�7�`�lX��1��Ƚ�))�(�K�g�kWΕH������o{ұ��!9N���Q��H�_�8���Kg�M4����Yg��k`�(�C�k����Ɨ�#tr���k�b/.T:r=o>>���ݏ�����7�կ�E�KˣQ,��$Y8�g6��&�d��l���&t\�J���
�����v�H�,`�4�z��z�D�rR���vUt�r.�����$3G=8�v�V����<��f�;*�a��'i^�ě�Wk�K_<�;�o����i�m#��#GL􌱣a��z��[��,m�J�1e��7'&�]hgW��W�7L��tH#���y��}c�ks���d(�h�9\�>��`d�-���(�T�N؍�85r���Z��s��g��&�8���M��|�S�g<�����~�lϦ�G_������hr��D}�g�ժ�{�֤�':�����d����<��5�h����
LB#�eKr�����_�ﵡ����'F���R�{��O*l��˪,�M��xk\�t�iM�McT�:��Tt��5s��1�`�K|�	67~��[Yu�wĴu��
��zcu��kx�6�2n��f���lB��a�(]kXٱr�-��J�<𗬩
�`�S�i�|�x�7V�v�Ϟ/	�	�N�=t>6Wg�8�|E�=��)Ctջ]ٿJk�Ci^S�{$�Ao�:�[�9$�!'q|k�G'�r��;�d�w�;�|ۮ�]�x�]�h���T�w�&�
�s��]I�8�,���W\�a��J9c��BR�Y�j��ۍ��f�f��$����\����M!��lW(5�3��Eo���
�V�p?�����uPt�@��C��x�)���ucz���)ν���z���%�6˽�N��;?Z6!����skR�k�$��
�ÛN�X����Gۣ����ʰ���$*�F]{>j��X���q[��7�Q*_$˞t�ݚ#m!�a����!�vǿ.1�8�s��^�C\�oŷ<�G=]ΑPz;���۞y$v��v�Np�g�뺷����~�~k�f��;��g�8��Qu��s�JtrϠ�eE߉�<��~\�;�����M%�v�a�
�㞼sQӛ�s�+�o�}{�p�7�J��� �r"6��q����.5tT���5眝ϢHg�F�l���1�6�7�A��%Unj�)k;�G5�/]:��,RvNB&�v�L�w߮|������V���.��r�>Ylce�-�w� �v�Z_>9�)�ˤ�������K��a�$01��
soʧ"�`ęc	J6
*�E��5%&A�C3*#l
H"��JLD#��!*�%�%XB@$HFP�aa�BD!eBX�3�}�]�Ϸ����o��lvEmE��}~C?������މľ1}���:7��*K�V�[t˘�/�,��E����.us��>V�m������¢%���O}�%�����q<���{_<n�bz���NK���i''V��5����{K�zhaT�b�}�����Ig3����zy_�j�>yu9�s�s��y�~n�<��߿[W�:�\��u���kl�ƛ^�oY��z����[m�=0����<�����z��C��~I罻r�~�Li����۾�m{�qo�]�u��Ҵ{�v�g��4��痊y�~�#���{ͯ����Y�SO$;Z�1}�w|�U[��w��}�zq]|m�Yg�]|w�^�s���r��\:�/XR�xC^^/�22F�=y�v���UXt^�����4���݊�t�]�1m��E�[��q:�������?ܟA��Ia,=0��X `�U�Owy�_;|9���~T{K�~����k��Ph����38�s�@:UM,�iNr�P�j�IG<@I�o_�m�yӎ8n������ӯOy����d�gΞ�	��9�R��8��on��߱�R-��������A-=g�Ǎ|��]1�ݸo�n���'���+���A���w_}�g'�F�{�ԇ{�k��yb=��o��L8�_^w�e�ݲ��W�};s���*�r���O|�w�Q6���[����Νz�q݋}G�q��/kz��Xߌŝ
�:��g�g�;���9y�nY�����b����'蓶�����aڝ�^c켵��������(i�馃�����A>��a�۝+xzzs�]�ͽ������7��{Y��-�s���O��7�5���>{N�ZF>�}<b[J�H9\�zeXu�ߓn�����ӛ����(?�U�w��b�aN�'~��{��2�N���HF^zPgʾ����ze�8�>�y�&hv��T��,�'?K[����s߬�]�㎞��o��^3�G��~ܗC�=��<�8���� ��8f׀}�i�AZ@|V(J� ŭ�~q��C��G 2Z�-�S{��d�H�T�T���S*����N8�R�Vp3�(�4."2ƶ����1
��l-X�貪�G���Z�"�3��:M��Y�Qs!�\M�n6�3D���ٖm�(M�!�� ɴ���o����|[�^�f�#���F�k�(i��g�������}�]}��<��JW�5�}��9z[�F��9���8�ܓ:;��ZzA����'�~�Ҝz������mk�����~a�d�ǌ�"mc���F6RA�d��z�F)%M�RIR��vr��:�c�����|��׿�E8��t���/���rv^��d���<�4i��˗��ۅ���Zz�:�+^~>?�j)ѝ=Z�~�S_�:���8����U����/ǩ�M7NbU`����8�p��i��4;3�������گL{t{e�k��a��Ԏޟ&�j_Lo�����ϝ��BT�װ�#�)�$�_H5 ,�[p����ڏ#�A,4���T�4l���6�*��q������YD�Ji��,ȓ��3��$�0�<_y;��?�����\VmU$M�7�ﹾ;�䱷��f#��|h��7����L��x���ƅ���L���2����Ǣ<u���QMW=�/M2��M��r
9���mt�|fU��Q5�rr֍|d�(12}��u"�<0��OQQ �@:E�q�:�CL82��:,e ���H��i�94�OZ��XH�m��\�Z�[R
eAO,��(8�0�,-!UH:��QJ����#���h���_��K�*����0"�D�4����aQ:�B4�4;	��9l�<�M��8�q(L.�,S0���G4i.>�Y���!R\��M!�a�����1���ݻ~^�׬c��߬4����o��8�7��(Y=�/u�}�R�a���M�	Ȣ�E�1�I�T�����jM��0!S�!%FvS��BR6VYM�EΡi��9�@�@C�ɵMeG!MA�	�D�8vp��9��(}w�����X�RZ32c��͛d��E`E�E2�KiJ<Qc�!TT#q�!�����	��KA�%H� �.\���ǇC����#=xU���DP�:	 �- �:h�R������vY�Ny0�I�dI���B�E/˩<��T�H%X���t��μ���M!�y����S�_��]N��>�/-���ܡ�C;�`�G�{� � �� 	P� �d�eR$FP� Dww� ����p�W��_"�yp�a"�;��Jr;����#�`r	���b���{Q+�	r%�0��;����SM.����U��Щ�Xq�(�5�(59%ǎ�PA�a�T$%� �>7�\P-�
����gJ�iZ'�.YDz�8ʀ"(�XΉaτmk��bDB�M�1Ƣ���B1q��ˡ	t�m(���$P`�H��U���N��<�C@塋\��B��$дrH[G��U�L֦zI�X�)��P@�!wV��VtR�2�^)� �@
b�d���m�SK�L����W��X���&�cL�0[F�uLj�KW	
	�E��z�Faîi�4a�x ���8�_�6aʞ��$�A�
�]0���Gc�m��V%!e���8�,8������%#TE�Lo4`�$�#�3��I�7`p���\��{��D��U�`R�Qh�!��08m��!(YL�X��]i��\�H��>]�)�=(�2��BɮR+W's�P ��kg\J��	Z��Q0�eA��y�"��V����"U� 1�g"{ܮ/��A
]�38�Bq��`2�`1��EBB��O&*a$&�:� ��a�����B�P4����q���|�)��]Z/!sUY�BHcI*�vX�D�4zϙ"TkF�H�9BCK�q2��#�y15b*a�k+^�nGl��$
"�`I4S���]J�	DU���#�J�@�󎲈�U*HH�Ү	FX���� l�$�}C�E�4�}�um�[��wNo����r=k��������M�o*�2�B����������;��^��~O���K��7���������x��s����znCs�������y���R~O�L�>!_g�r������w��+C����o����G��)�ߢ�X�jT%&��������D'�2Wձ������k������������t����;�)�~��Y�o���W���/!�~�&�{��y��|��j.�<_ �ˈ��'����6�9�iR��è�|S�w���A�ya�B?/!�y��������6�w��G	A���*������W�h\��oC�m����7(ȩ伷�xԺB������?��G�e��|�7�H]���2)������p�{�e^Z�F�M���V��~W/��lo��Cg����~g�-����y?��K��(���W.:�,M�7G�L/Q����y_/輧����x���ϑ��q���rۿ�4���������<����m��wx�"��8�?5��`'�����=?�Y�|f�=d��z���Ǭ�OS��ܓ/S�yo4���ctw������y�k <��)��
~a�����xz��H��r�_o��5u����n����Wg9��� yxEiR!P |����'څ�~���h�S��]�Y��<?|?��g���*g���Ĝ���o���}�l�q�(se���3���C����c��
PQH��h���Dǳ�&��^����AY�<�~�ߎKU@B�8~;_�)���f����"X���!,�M�֓l�D�9s�)s0���L�4�����jM��50��c�א�.,< i��G��î]�ml*���4ǎLs+�N@�8����ԴX�VS�FS�ʕ�F2�T�8C�+3T�FԬ,Fvm.,cڎGʈ�g�9@hHИgŅ�řbN|3Ip�~	T�3K�.r���Aa��m��3����t���L�� �k�,P#��d���6M���%��6��],E�r�&�ۡHȅ2�8�ZT�62�+0����YX���Z*�;�Аxe waA,��é��!}�[���aC��K�"
��d�PƲ�-�q���	�{�HP�5���%ae�x����'M�A�V.�u\`Ƭ�d� 1j�X��,R^e��r���b�r�]#�9���CD8�MH@z�8Z�����ؘ�:���qp����tK��Ӭ�$��3,��͖	���9�,S��B�$b��KE�Kgji��ՎImh��J5��$��V�1� x�o�-Ӏ�Dh���L��	�"�b�Y����2Ċ8&eC��1K�r��jZ�DD��jb��$�!Z"u�V���,�A�ԋ�xB,,qJ���8�Y`X�>�A��Jfj�N2$2���|uo+A��w�xHKP�l^b��܆���L��#L����SzX3�\�ɯ5��r�k;t��7���ה�&j���M�']�_����|[[��G����<B� D���)Th):�9���S��X���^?�un'7�y��X��х҃������C,9�OI�6d�Č4����G�kE��I��l��O�c��P�O����),�[[�~Y��#$:k�C�[���d`t6԰F��Kl|�����1�6���R"噪\�e p�eeM�4IR,�k��]⅋CR�p���6��Rᥟp製�6�$RM�`QY�(��E����sR�mZ��z�|;)L�]B�\OS�>WϢ7_usV+b����`�D��G��ܓ"��̽7$���â�d@r����:�G�Ҳ�5MX݌�RQ�H��Fmj�?����sj�j���u�LbLű���$��Ie�� 8�e'!F�h1�� m�cb#4XЍ���O��/X� {!ס���Ԇv �˱��@\N���:v���0�#t�ɣa���d�ƺ8��[REZ��X�i�B���9ub��µ�J;�F����ӌb�!�:%	����'n�޽B��bi*6*{T.um@�	�lS= y%�(�a�2͉9J�;,!�Q�Ӝw*�cZ�b摱���.n�i7Q+�D$��NR,�%;�9ԉ�+V��{��ۦؤ�/fj����f��i-��^b�8A���6�6�1�
�Vހ��ҁ��r�64E�~̴e�ۄ�!h�ٕ94�
Y|���.������k@ʓ#�������P#�.1�M��z㯭&��h�rU�ZDI3BTFK%�N3$]��:ޤNhð��R�k��@r�1CȒW�(gFV"F}k�X�O����������ym)b�*6���fX�����*�̦�h�cfZтX5����+I���R%,*�a�
�I�|����GM2��T ?��#�3 �TĢ�0�[L� �%BB��!��L�@���i0"�pbA
##"�ZV�
PU� �
���9 �i4�s]�2)IV�V(�e��Z�j�@��ZP\@�T��LJ�q	H��)Tq"�Ҫ �@�1�\H!CBD*� Ģ H@�!\H�J�! JQ���U
UZDq�
��P�RR ��4-
�b�P
q(� T*�(Ы@�-����E��TUnmrܴm�b���A�mʍF��5��%Q`�t5F��b+��02�Y X�R%��Jс-AX�#�
,H� ��Q���d��;<����Ą��#"$X�5E�,X�6�QX�DjC��;v1�(�5�Q�UFجm���	�͹�i"5	��Z"�j6
�h4ZL���4mcZ*1�����6���wub,E��E��lX����b��cZ5�@j��ZM%�Q؍��mF�Eo���e�/�g�3�����c���������H}������g�>�����>iO+�^�_��ޣ���������}��#��'�����ܻ����>'���s����/�}ߓ{�������~��x�Y6�������o���1�_���>���g���_�}�����{�?��?}�>{����K��'�_��ڇ������?��=�|ϵ�|����Ϙ�o�?���������_g��?��տ��W��_���.���J��֍(XFF�M5Z`�X�I�1I�d �j(Ʊ�!�cmE���T��F�Q�MUZ�V�h�l����4lZ-��Rm�lkI��m�j�ډ,�,l������m�hE�6��kX�Z��2Ȕ�R)J�-6-F�֢��E�Ņ)b�hE(U)A
E@JH�R�Q)J)B�T�DH��A�(iQQh(P
�iB���)6ִlZ1����QT	QlkD*A�1Q��F�VE#�"�&�$F�P�&12�DS@F�ͬ[Dk6����-QQ�*�l
��@�B�("%���lUckZ�UF) Zh)E���)(T�i�F�JUJJi� �V6�
ڍZ���`j��Zh@�P�TiV�E�Z�ZA�QB�(R�P��ڊڍQUE��h�kb�*�-�j6�+E�kEj(�JZZ�*��E$�DUO.a@���lJ����!	(���_o�8^?�{�Q���� /.���}?��?��{j~?/�>Y����6����<��~�����������k��~g����_��������x�����[���������w�����>g?��?���'�o�?�}O��������[����˟|������?+��K�>f?��~7י�^IO��xv���)����������0z�~_�����?��r~��X?����ya�����9���0������7x��S�?����=���O��z�?٦��<'%�����^���/�>�!�=����S�>w��N��y��%^[UڛT�*l�G�����[�T��"��LH����,H�$��D@4�I2�����J$lI$�ɔ�1$L�!)&SA���C&��c �hҒ$�Ƒ1��#`LQ�DF�B"X0&���Fd`1�H FDBF�fɁ3Rj`İ��I(�!��LF��"�	3J
#��H�-�H���3	D�HLȑ(�21�S�!$j1$���LAI"FF3PDQ����"4�M0h��I�1�B��0Q�#��`���$bE(̑14h� !��%!�*i	K"Bb$Q3!&I"�����&�(�I�$R�4F�&R�I�B� �33 ٓLRh�l�I�)6Q(�A��LȂ�2�f�f30"!�"�d�C �	� ��f������	�&i"�6&`�D�h1��`�
! E��f�D� TCBi�BH�#&Jd%!�H��`i)��1 )�&	 �hf�Rb��bQbH��21�ى�i`Py�T�0��T|D��L�<�����&�����������?��k����S�����~��o�����/����?g�c��L�M����������?��������>��{�{��?��?������u���|�|�}��t?w���)�?s��_���������~���'��g��ʏi�1>C�J�*:�xIPL�L� ?�@	�ZV�i 3�*�p�P�x�P\J� R�i#���
EvJ�*��¢y`4�C � ��!�
P�C(P33� F�W��IT2�*�"1��0J�DO*.�H�P�!"�^G��;?s�>7��?{������[�}�S�*7�<�t��������t��s�=o�������?���W?��`�i}W�G�������[�>��]�?��������K��=��w��|?�����/l���O��O�����:��_������������~H��� ��_������������I�^���������h�_Bľ�ӫ�_a�
^���/�n�a���l
�������_�d�^�࿔�E��vDT�:\���j+��h�=h���dIU�B�.�U��H"���rŝ-��y2h(1R@��\tV�v��GT�|4���0}�_�����l�R��"	ĝ�K#�s�Y2�MEV����*�����Q����,�2�r��q^�/��]�����3#t�c�}��7�|'6 ��l9�*;9ͣ�B��˜~CDW욡� �W#yf��8İ�'aj�m��Y�xx߆p>� �`6�,�f*h�p ���nX(�$}��=�(��{���)j$�IRE���T�z<e^ �#i��A��.� 1:���Y|Q�=kv��Q�O�w[LR!�4��z}� N��ȝcZ�i����Ǳ��� �C9��q�8D��;NI�$���C���+[8�c���I�a׆�p�Bd�[Gf����$۶�ѵp=�������5�k�h�#�R��z�PD�X[U���Z�\�y�p�F�h�ղ(E-��̩EA�UM�3��ƅQ\;4IF)�%"���U��3!�A��Z�4s��x�#�(��L���p�b��Sj؍��d���v���[q#(g]e��^b+@�qPX����I/-Za^4���[�a5�MAD�����xŔ`il'Ҝǆ=��v	���p�FV�#r|7� ��9<1ػ�tɤ��j�!4�E��[Nc��I���/WwOb[8n�r�]� �Uգ=�Yx��U��#f��ʔ1 ��_�AW�Q��� �70J揢�s�l��j{Y[�շ��iA,��Kڀ%`]�%�D�q<���MGlF�	p�s�u���b���!�QU�[���D`C5-�}�w� l��u[3�;���wu�0���t4\� $�
,�(=� �"���'�c~c�ӝ�:@Ҧ%�Į��&PiڌR�1�Ƽ*:I�V4�HJJD�t�H���Gv�BJ�V�#����6l�����d!����@2�
#� I��%&��ƛ0����� b5j�!
2���K�(����	�Z���>x,�$�c$�a>��L�e07�̲mI�m�<;P���r�<�vpf|$�&Ri<L�I���,�ę�:�HL�� ���;#^��Dٍ��v�K��O�ϩ&`g��$�|3��갢d�<_���3�$�3O8��)�[�n[ݾ�͹k�>���U�C��l�;x��pg��kf2��L�o���LL����'}Y8��M� #��.c�C��%�0�������k ��ک��1�|ff�NRd	I�><�$�@�g�S�����`AP� i }"�He �4( 9@�"�)W��A�p �R�;R"҂ i*�J�~@C�����J*�Ҡ��@Nr@ސKf܌m�2N0 ѷ���0�a����L_�&٨���4�8p'!p�(S8N>G.K%)�"dӉ�&L�96����������>�6N��l��K^�6�;R���T�[x��i [0ꕣk< j��$1��MP@`�5�q�(P٫H.�jMR�J�I���gUҚB�]�!�	��vc	G�)��8�02wђ<���'���3�&�4�L�(d�Y��-��Mq�LB8����K�MrbBgK��%q#��tمMPk�s�'(�:��M%1�^ k����s�V�	�q.�H�[fY;p�p��]�SI6�@�����8r�(Ļ����y !8H d�W��(+$�k6*0� I�����������������������������������;���ml�j� 2 ��@l   (�
.                        �               �(  ( U      :�             C�T                  ڊ8� �  
 Ɂ���`     ` @p   `:4  AB  � 
AB��(��      /`   3�`      @  ��     '0 ��      �%u�  �      �ERT/v�    7�      �)X`P     � \                                                                   �w�       `       � B W���tHP                                  ( �R�   @   P                  @  	�  �T��jUޜ���  z� H    �(  �|   @ � �U$PD HQ@  `   �   (   tO�hJ� 8    �hEU?�      &@T�'�A�b'�ɠTi�=dɧ�{T��j6Q�=���eOԞ�F�==M���62�4����54����  �A	=mM��� �=M�ީ��z'���ښ � =@� ���       4S�	UTɨ                              j~D�R��00` 0	��� ` 01&	� `   F�CL `$�IIJeF�@ �=@�M Ѡh�4h���    � �h  �   �  B�$�	�Dژd�dhL�	���&������� ��i�i<�2bjcF��z4d�=�~�S�F&## C�MOI���3J� ��
?�@�0!`�I�X�h�y,�!����'�t��)��g��}3��Ć��&��\>�UD�� FO�����k�O*e~O����F0�����f.f͖���5�h!�D� ryJ��C��n=M�N9�/9���V���B$�C�pcǭ���a�I�����
��-���8ӓ���s���l��B/������}�ĳ��o�,������� B��!w��kHVn����F���M4Ά,زd��Ix@x	f! B�����V��T7_%R�`W�����ǹꧪLV�A7�~=�$�8�A�P%xN�wf�&g9�5c%���&-'6�5�qo!��q�����b� ː�'QV`쪹���.5M,YХ�,���(�B��#�^�b����~ڶM�TI�����DM��P�4Xn�8���N��'!T��wf��9yovmy�{������* 
TN�7��V�����f����Sn��lng�G�%fE"0�x@LT-�,3��)�d��`���6I�
�m�)/����}�p��!׿;+:ܱ�gT<~�e��j~֌܎�e�a�uq��\���̸��׼����x���$�:\)xt�~�k�i3{C�b
�ѧ}f�G��G�������uW:�,<s�O��9��zA@�eO��3ڱȕ�:M|�F�]L/N�m�~��s��C�Uy�ᡸ���H}����x�S���1�*�����N�8�ԝ��5��el�y-���4Q��� _2@�tz��j%k[�O��wLZ�湘�0D��U�I�%��L���Fd�;��WN�ᓡI^$�;B�h�k��a�?�ZY�OS���yʫ"vy��Sg��+>xM�u��LS�+\��/�#Z�c���L���F��"u��A����
I�X���[7�:ol�[eϊD�S�����>m�B�m�@F%Ć�L�1�_��.�JKKꅞ�I��[*�wF���6�E��:Q�N�nѣ<�c�V���Ol݊qo�W�Q�u{^:�Z����jݒ6]΋VZ����1(���i���e'z�WT.��&_������d� ߦ�f��$��f�YM�=�"D�6l�{B�Є?@���R���ԍ�|!`�Wf���t��[�+; �7e�������<��cMx�q�""8n6a�h�"I��a  �q��(_c� ҂%�E�VX�����{5�j�D��"����U"gU�sm��ۈ���;9N�v$D��J$PJ[O�ɷ5۳w�q&���bq��Ea��DX1�q�5cK���ŷ�SGi�{�'r����9�c��[�
�ϑ����!�y9��-�v ���?���σ� �/�"��|���Ɉ$�A��AUD?���������|t�GΞc��g��ea�s,
�	a� �:�f���/e�fEΗ�n�Hy�jN�03Kb�i�ȃH���KO2���q#�Z�gX\,ɇ�!�κ���Ey��v��x���d����� �K�g��X�F�1c1� ���1��"�M��/���c�HS�R��[V[Y6߇k:p�ё��S�`��W�,DI\]������<�HD�� BB�����:��(��y�f�y�$��b֐�Y�IN�s����"G�!d�PA�Z�� ����j�o�
y((IĢ���0� �����CH@B�Q̨H�f1
-(�Т�q&$TS����SIA@)Q� .�����Z	I;�n�	�RA@8Tp	lh�4��?qm�cI����	M-5��!�
���_E��u�TĠ�~YA�	aR �Fe�ID FaF %FH��I	�}��Z�Pu��ECvEC;��9Z� �$J$ @�,��R� H�!*��J��A��x���Dh7�U��n�P�d �]쪮���N+����wa�A��U����x���w^���o�~���ϔ�oW�޳���k�|��zoa��|��y޻�9~{�ﾳ��λ���>����/��ޛ�{o���ˬ���~����[��UaD��"�{om�����=�U�7�WY�����;ר�}����O��1����������������v޳�{����s|�O����[�w�+�=��y�W]��sӦ�*� �(��|��u��Whtp���ny�5�y�/]l���on\��˷��AQ�S�������n���M|�'T����t������)�J�v�n��/z����9ӡ��߾p�mN��Q�B h�q�N^��R�ch�/86q��r�N�L+���=�]���oqotq���;W".��(��t.��[�eKXm��<��E�HK��>��!@CɎ,l����?�q��J�x@@@BR�u�6p��W5��# !S��|���HBۻ��q]�(!?HHS�+�Ï��C���ˈ~��q*{�s��?�� B�I[��0���㟷�`!�{�  w�kjE=������G�9 B���;��#�� _�QC＾�i�:�W����W��>�!!  !ď���Zz��)�������B�� C���17(��J�H��kq   g�N��"��Qq�@B��G]�!����� ��_�������|[��_o�D �!
_��C�Hd Ux���<-����guUW��Q�n󭂪�[��o��@B	�!   �i�	{�_��R/�O��!  C�M;���i�w�g���_S��� B��w�~=����  !��|��p�O�ٗzWf��  
6z�Ǭ������7��pc���9��g���\!إYg@B_FU.~�O_������5�c#�,BZ<Gh�=�U�  �+�����}{�D�X��� B��|E���7_�C�V���  !V����8��ް�!����
�!���q��}�`1  �e9�ga<�Ć �(��+��F�=�  !�	�a;����2(�TZjv� �J=�N^���d���u����  !dF�a+�I@@B��"ƶa��ih/z��x@B�� $�1���tO����!=�_�XF�׋ )��9ⷌp�7���Q惯�� B�x>5�{}L@BQ2��c�uuH�^-Ѹ�I�V�F�  8m���3�5�׸�ݥE_9���W�5�-L������ F�m���#� ��Dx�=1��͚ŌV�T+a(�~+�(zz�,�c{��)�U|&,<5�L^g��8�!�A3B<Jks��$�א�@��� I!�VZ�UYl�*�$u�<Fڡ8����S�@�K`@�-,���ƿ�;5��)薩V�I�u��M_4k,$�!�A�p��],49�����+�i�^%۬kƙ�=эh@9i�.(;��5�':�[|������B>}B#F]{o66� �S��o��������d�B2�X�>�_F*I�T�h��ޞ��Ô��>+����fw��oV���,��J��tp����d&:��O~Lz}{�� ���_5	��|�<��'F!
�<��������E@!�5�ĩc��{Jl
63/�*���
��:u��Ft�������l�M���Ek�gwm/[�Sn���#ͬ䝝��N��S�m�a}׮�b(�<�����R��)/wkZ7Y��t��N=ldX��3������i��do�@ .-s��%�Ks���t�_j�Ouj�'�%�O@Ia)-uqX������ �>O
��� !&�Ձ�����x]|��,T�׮�R���!�jn��1P����,8��d�x��=���)&���(���b@�m��b{m��y�KT(@W�"o�u��a�!���)eu�꒑{�0�[��aҥ�'�$�U�#S��Cĩ�Z��2+�ȧ]Y[���
�Ut�vLL�A8LbX�b�,:�{���]q,&� �(ki�3CWiaIiV,K	���P�%�qQ.��$�F�N�-�ճ2�=��!��%ྥ�`�fJeI�_D�@�/�5���d��N%�j\[���z��l�q�_:��P<�D��5�[����xt�Ɯ�x��p��P�)]]͇�ճ�n�\݄�U=O66ˉ��д��mp8�ePZ��J4oY��O_�F=���J��r�@��>8J�.���gk��,{k����1J�[R4�n��'��;G�Ou|�Z�U�J|K�{Q=�U�
�����c��:$���P�`L/Z�r�K�;H��f�lvc��\��
���Ϡv�wP6ֳ<J��2�Iq�y_{s��Xp7in롱���^$��&�3h,�ϸ�
<k��*�x��D�Y5i*y�VZ�M3�)�#
cwz�%u�0�sH�JO�1�I}Xѕb�<{�����)��p��XηQ�=;2�1<�t,8���b�w�}�=��l~/9�YF�m{��:siF &[�a�Z08�Ԣ��y��㭧���
Z¥��{�W�h/�ô�_K�^1���"����[�[�DP���<�6�
F�$x�4=�8r ����_ 1#�"��>W�|5nޛ`���D��m)@	FJ�D�$Fa�.�F� ��wheN�_U��r]��aH1JK,ϒ=�Ѫq��18ƈ��xt!`��~�n��|H�ka��Ӥ6����b�<>�#(�iOդPQ7\���m�����l�1f�,���zZ�-�����,�@�Fwޞ�f�RƳ	��!:S���'K2:�q)E�����9��ж���\g��� h�|��J±�b���e���'�I;�(II)�/�{����M�N�$�Q �@��yZ��]�;U�9��zՕ��F0��7],S�RzZ�T��q��111  
V�a3���z�K������D�@������4pٯ�{[����f���u�Ő!�����1��Y�c���zɪU���x���a��^(Y�ϟ,�����DO A܆���"DXok�{���H�V�P)�ƫ��C/��j4�����D_�_����a��~m&���72�շ�`ӲJ1eb}})K%78�=qWik�J�z��-a���X��e��Dgn4��ēv�ڡI6f�xօ[-e�$9�a l��O&1���@G��1Ʃ9�
R��
��>@=����X
���@��)(�'�Rr͋b���q�k<��N�>9�#'�*�[_s)HJ��A�n)�DXg�'f�O=o��uOLv�yB�����{)Yv��$'@�|���i22.i�
f$8z��e΍�at�=������S�=Kn�����(��n¯0IN5-�BXMͺ� �԰Z�Rs=-�W�����a.�ֲ��'�{�Jxf��j�/��1���w��Y}Kn��:�_e�%���,&�}tQ�����ڒwlcv�:�������{Y���Ɣ�"�(�m�V"*��+�*��&����,r���H���P;�@	čiA��&���@���	,_"y�_!� gs��"$G��3��uOʤ#X���'��Bv�~g�6�U�(V�;�{YM!�D�^�zzt�^Rŋ�`j�����z(|�dOF����a�%>��R�+,��t������|?)�oI���➘kI@�Лw��zz~!�==5�xW�9��b@�,������i���[ض������K)Y�Դ��Y�i�[�qC�IF��D�4��{�e�@Aѩj���DBf� �+]c��d�J�o�f��8[^덭���\�$DS��M}����W�SŌ|K}[8�s:�+$z��1'��>}򡯓)K���!_8j�`m�\�!)#�c�1��{JqhYY��HB6u�|4��~9dOnaV�����q��D���m9��hXf�ʥP<Dfq��W��%��f=1)���z��P&��kE@�zR!!KVҕDǱ;��F	孈�����k|(�+'l���la��8�k˘�&2����*���H^��0�!�\g��v��Ʊ�<�k��
��QO`���F@��jY�e�N����Zl����
�=�ƾg1��fXzuq:t{\؎Xڤɬ-�S��7�+)(ZM	`x�Д��ј�n��f����͗�n�@�K�$�XF@�2�u�!���h�XEf)X�=� �k뙰�ik
և�ݤw64$���+9J�����9Yք�ӧu�y�<B�(%�o��YuM9������Ж��jv��r%���uvi�`<z������9{��x��HB�%U�g��u��ҁb�bL�@/XZBA'BZs/��Ɲ�����&�6_5�6bOoɯ��ŀ����bR5c9l#5q^z,B�W�@���'i�Lz�J��dy�iH�wK!����)�Sݟc���!u�[O<���^�w��~��}IC9dH6ЂF�4֥|/��s�X��S"�_>=O����B����K�%��w=�J�{&���|�W�$���f<L@�g`1�e�Oժ�xI���#���3L�n�U� ��(��HKX���SДs)	�]-�%z�ކ|��S��8�	�,��}D�j���ʒ>�(�Q�f˯�HAe���B�����Mu���6��N��IX0�����be/VU���kO A��~q	+=g=/6q��qX�;��I���|�7�l�/k�ο�l�=�1�����s��~��:�1��G���?������[�������%�b�Y��_��?�����'��j4�3�x������	���`��?�?�g�`S���ZPV?���]�+/�d �����e�����;K�"'���=����ݑ�=hG�F�>���{�/l�/����s���H����%��e/�#��y���K�?���{�`�[��_����y��/�*w�!��L�ۑ'�g	�QmW�hfӵ1�T%���7j> d�W���׌�@]j$���+_�z�{ɺ�T�u%~��J�~���-�z���JC��/�#䑒R�Y�����������K�O@	?]c, ��;(e��I*����.$N�%�"$H�A�lq.J�v�İ�洒�i
(L��*�m1		����aq����D�:^�%!8h{U#9��<>�&���Uy�ؾN���|�,{�����)�#T�*Km-@��vak�If=a,�]�NY^-b��m���]{��Ht�JD�`�˔��y��S�U�(�)�M׉��7n&���qբN`[�N�iYM�Ma*�i:�N��	:�h2/���۠�j�f.�ӹ�p�z4�3�䡘6�='�����T���G�$�M��K�_a|���mf,�4�Fwk�/�&0��K.$,3���,a�T!ζ6K	&P�HXu��eIl����e��8�[��!X�h7؝��9��X�@�g��=�$H��Ҕ���m۷{�f�c+#� DLz�f%�%8p���/��:gЄĵ����ϱνc�2Mc����J���-a����XN����ڐ��D�F�,��&|�YH�,�� $&"LH��g���eD�T8D��z���B|B��y�!�&��_Yxk:�;Y�Lh�g,Ё���Z7�{l<K�beP��j˵9��N^��U<DH�e��<^ҥ'	��r�Ù3�5��ѧ�H�c.���!�9H��TR(�^b{����QE)YIJ��2�,r�0=)�Aba��'�Z��hD�� �y��6/B7ϸ�8�2�0���|��DЋǬ�8��D��2��%�9��J�����Fp²�C� :Tg>aW�N���K۷Lt�,ݴ�͜u�k{>;�X�8�U&=r��A�\N�n�'�	z�o5�=��d�:�bSҭ����u�"9O��^�HV,��H��m&Y2�s,(-�H����[[���;t�k�:>�۝���v n�� fЬ@�Y�ɪ�<�Q���jxb�Q_���)R*@uv�R��|B"��K���v�0}�c�2��@	��H��:�Y�(1�x�aXJ��Kh�:ٟY�K�[� ���U��{V��HR��3>dD� ����Ĥ�:a��bZc�T^da,"�� E`[��v,<�T���z �ͭt(y$s�R�����z�[Ya��+$Lms/����Q/�R_R���@�� Q%Y $ �"�G�e8r��@�v+|�+IC�H�U)K3BH��AgE�=�B0�Q�k�z��p�,�Z!�|���J�0ENm�1{>��# �|ʑ!8H�|3�#�@�'$b� !X��� �,�>��`�0�>
��� B�"+耑A���BQ�X�8;N.丰��N�gA�b�q���(JF =f2p�۴�y5d�$���mH`��1ҍ�S��d� BB,����U$	"���XT���R�(*ZK��������۴ն�� !��d :[Q  ��!*��R�x^v:ʹ��xA#&,�ζŊ���j�f��Ҩ>���8��� @!�k����z�BE������em��b�a������υ���Ҟ��<�񉕈�X{Y-�e���K��dkC��w������\6��)K��3��z�x�R����ڒ�洐-bV0 ����B�z���Oz�� {�$�:���%.� MA�JD!��V����D��&L�)	~�T�����3X@"���(�c� ��K�׬�p���		�y�M�	�*2N��s�;X�R��G<Q��k�q������E����Q;Ǆmh�C�S,X�0��^��d��v}}�C�Ss7��\yX�  ��xet�K	H���v��ݻϸz>ձ�z�$ /�J�d�)5�xS�`�T��$ORB^%�s,�^���B���cP�a 
ǙIk�` �)kϏ	(��)-��LIg:�$���� rÔ��ϯ������O���͔S��8���+ݬ�J���I�ޚ%�.��"!�N&��3觐H�����&��,	���9��%=�,����{��:�������D�_q=� ����ܾ��F���/X�L�u�!8���bJD�=E�f	���=�;���)1aQb.�m��k�W��Jz�1%_ q�q�y�x���V>�����W;5U��{��]��^��v���v��{r��,OC[�[Jc��"(� �X*B�f=1�s6�>�����X�q9�b�DOi���q,���i�����ľ$FZ� r}.y!����Ss��z>�9����'��O��Luh=��f���"�=h�=�gwK�y��h��ow��B�2)�a衋�@���j3 �	���[l�&�!	ٛ:�r��[Ͼ�ބ�RLKl��8�kg.�wYa��\��-i;1�l�xN<[J<9Pg�s8���ZR��W�񥔪'�Kc()��Q��) y<���(y�N-���IQ	���VGY�w6�ԍ6�����E��q�LH��YOx��KQ##<J���L�#�$���@��X1��H�̲��m�lz�}�А�� 38���}1J0��<.���=�{�eM{���i����B^��Y��5HNt!ZJP�ǜ� �.���g4qW#H	��|��#ݤ��f5�+�����b�m�'��a	㵗3�ډ���.i���_-$�VMRc<n�L>!���C�VԤ$'[bYj>_0'(L�8�&���z�7��S�	K|!:ҞN���VW�3'����h"�P@�L
Xk-��%���
A��Zq�1x�H����ȅ���e���)I�ڒ���πќ^7%�'eHŏ�-f�1Ω  V)ka�eB��:�]�ӻ�# v�
����F>�5O �u;�L��y�.�#��vn)(0m-%ia+�o�^�0z�e���x��*��bLB� W����b��t׻^���	���-Z��%�[��T���SM�P����,�ŵݰc=ێ�lb�����#������(�=�"\5_	7N{,�𔧪�ď����5�����'��Kl-���i��؄2��Kkz�#���挌ݴ&�K[>����N��PԁgkPc� � �����}`S�|�S�`�LN�C7į+^���m�_$"��d �N|��$B4d�Ǟu�6��#;��o(�ڄ�cu����\�t��	z-� �����"�B��i}i�K��w3OIa$"����� 8�I��=κ��O,W{)��c��[`�bXTl$I`E�2��U`�@&���˙�YMH��Ʃ���0��N�ʲ�ƣ M1�.Y1��[�F
�
�8��m��K�y�l�"G)�!���=X�q,=V�ķ�/��;p�iI x̌X�kX�L�o*�R��Vm����Ъ ��62 yY��d��Ϭ""�=�bq�IO;��"|~z���!<Wh�o�� HN#������_V$-�����0z%$
|����2�)-�!_s��ղՋ.��C�1<����<y�6�^E�Fq�&j�1��!ُ���3�c�*B���8yӊx,"�����{ֱ�W����)�F|�')�׷v�!9g/�����.�ԙ��׈���a��.�ة1|�7�	��X����<nq3���������<3��U�$��)��<3�y����
�xG�˵o��D��\T���Sˮ%��E�V0X�q�Vl��#���x�K�t&�_n����%��>�_Pk'v�y8��G�֒�"IH��{�y=4#��<y�%�|������Df�k���΂�cW��{��A-(�� 8�U�0��������a$����|��������C���w�p_�����p�c��'�i���?�����RO�GG�'I����I�����?���q�7��LT��@��H�g���߽�\ϻ��?���-��z�{������|?��DC�
]��P��Ԃ}G����tE ǁ4�)������5"�����h��E��?�A4�B���'j�˥�Jmv��q�~م��o&�3Ŭ�h�3^� hj�F�d[�c��N2G�"xz� �  �   �E�@)��y������&:�oQ����Γ���N�����"�4q�uꎭ�_OSMv�<Ū�,h�3兓u�E�|@��^�8���L	��DM��,z���i,^�^��1V�"��31�fO+�.Z��QUmU�_��.�o�~������-��
Ƶ��(R`v,W�P��iL��-W�ޛȪ�-&+��R�<we�F!"ҙ��)�5�vXd��ڨe��vBq��.4�P�_��b��ÒZ�Y �چ�s�X�<����'�Q:�<�E��������\~Z�~���_v�X�[�0���e��Mi42�I��x�.8��/j�/��́J}E��{����G�3��k�MOڽi�0,#��A���i	�M�FoN�����v�|�X�5fҞU��,ʭ=<Y�A��Ў�P��+��a8:a�.o�l��b�Ue;�Od�:@}B|����� ��=g��s�v��<I�M7֐�$B^׍�,�g�h�F�I�)E5�U���a���J�����#��E�ﲜ�T��{��Z"����u���t��'%�AV��'��#Y�����p3J���a�Գ�T\0��R32z�jPs����ťq�i��"�<�A�^�*�v�6c7��ZIx@RI�1%3R�5�k��ʹ,�
���JC�
U]�yR{�Óܡ5��5�R.T]��f�*o�em8M�ى�?rΫ5(�=�&\���Ź���h�}���a�l��0�zј�Sa�t�U@��8��Jo4,Y�N��Z;{&�IǮ�ˏ�<����Ӯ��;���YK�-�h�8��O�S�W�󫥛\�4��%8�Y#�jj$��HH cJAfC`�y�0:bdc�\���hꒂ91���YS����l�ѧL��LȬ�&/+�j��7F}��`�Bά׉Wk;��(��i�h�.��u��Cc8������#�o�t�\[�o8��i�I� ��ڳ>a)�W��V*o����� 3Tx�0�1ԕ��w��9�p��P�Å%��]�>�D\��ot[l��H�u��<����M�ۚa/�e�̏6=�����O�6�LZ���U|�:��5T-'���k�S� ;A<:�z��?4��b5%�o^�՘�,���aD�8�0�2s�嘄�F;]/{sST��t%]�S��Ė;q&�Q���a�]�
��<�_R1[H[�D�\������2)j�Aqh�%J�P>��<��+��6%G��5i�Z��c��j���z}	NY���4cM��\��(0dGI�B�x�ŪJ��OΔmvօ��P����G6�z�%1�g+�^h����N
p���E�S���+�# v���4��k#��u��V�¤�D0���)~My���!�6y�^�ь!P�R4KN$Z_|���b�_+ME������ǰ�r#�48��`]s����D��i/+b
������M����8z��o�PA���T<@�f%T�	�q� !I���ʈ��P�4��s .P	@�g����?�����������,�������'�{���-����������;�������}���!?�����} ����ʏ��m����H�o8���b_�JO��\�����D>���-�I���ŉ�j,���w�N{>��	���)�\��g��� cZ[��b
 /��+ eů\�_�m[�l���1vE��!ơ�9���+��J����YHD@y%�4zR��W�?�O�7�n�?��&�U�,U�EW��if#���T5���Ycg&-f��<^�Ƽ���n<h��}=I���!u̚�iα�Y�8.e��Џi�}"bP��X�&���-������"���Cp8�=B��Ӹ��9t����-��*��J�Y�Qa/%��&��U݊7�s��+nD�����&�^`ÂN�z�13�-p�Z|�z����荢.���j�ĝ�j1����6�W���� ņ��?٤�s~�'�ec�����<B8���[����4;�F�j�9C��8	��Ȩ��36�X�!�Μ�tQF�nv����֒O����@�@⒲�P8���l������+oK��D��
 G�y�����=�*�T�(G�b�z',�D�D��Z�>����Vk�.5*õ�!��u5^b�pcQ�T�����=��%<�`0���� �t��Hl8�q 1���#��N���T�A�[I ZX��܁��O$�Qz��!"@�bRz�H)���F�V�3���S��X��Ì r�����[�+�S�r��!�*��+,��e{쇱���0���R�>!�a�=�S��d�|���̬V�&�w>/�k��K�fLR|����U\�s�%~�x�x<K�t߂�sQg�Ѧ�X��n��{��i�-c/t7$^���W9/�:5��W��LQ��_C�8��t%�$1��;Q�bZq�^�cX����+	r�Ṋ�E�zcC��h�xɻ�*�R��؍�e jA^�쯭��B�`�NI��GseK7�2������UbN)�L+�g＇���"݉��/�sJ�<��ڨ��$�B��`k�7��;��E7��]M(3^�:�7���4�Ņ�S|�&���S��#W�iGJe�<g���Z��IT�,0 E�5�䱸5B[�R�Vһ��T�QǨ�.�gGeS��8!+��A.����6�0(6�g�Mh�R@�Ú+��bJZQI��ǅwNd*�֊&�~�m��
',�PQ�_� <tW�Z���D)�"؀�D:�I��
�C��2K' $��_�웞E�r@Q͋C�}��P���lT�0���K۫~[�O���=�M4�:�(�Ι]��*�x)(�邬�_�� �A�R��<J��c��i��5�C� �[ŧ��L���S㾖�I�~�mع�M�\��f�JQ��K����:�\���P�D��vL>�e��r*��֚Z�
Gqk�=�]8%I�mJF�b'cL�O�ӊm�N��B�B2c%�%)�I���V �-�p�1�>�v\L���ܜRx��L{�1Ж�ODA���,t��,�k>*�Q�6�]�NQ ���;
�L[%�C"̴b�*�^�4�$Z�	�����s�����`M��&�K؝�Ɋ=��F \�K���8�|.�2j�P2t�ɨ�o�7��s�m����VD�jE�.�n�ݞ�2w��H�*\�A"x�r�N�Ҥ�i'���=���s�~Q�E�H�'���"�i�e-۬,ԏy2$��iA����+�o5�oG
	�Bg���iE$�d���c�F� |�@�\��t��2�^�qs���6G��n�P��T&����:��!��	�����QcUH|w�>��:�����XO&��d��G�g�BӘwTb��X?Ь�P��>�+�k� {)��^<�^2��ֺ�eT,ozXn�N� ��i`L`������5��_~�j<���h�N3�f�f�6���(W� �X�(:���H�+Փ��J��Heq?���g��og�~,%�����F�+L�Mu�(l%�:��POK�%U�eXf�iTZUwI��
�g���Wg�6|��l��������T��|ӛN�ln4Ca��ݫC���
���۹��S9|c���\�%ۀ�u��!��T�=Գ��h�i�6w�_�f�@�4�}$}")�z�*���c�G���'��S18m� �r�!�	�hO[zUS���eB%,�Pt��%�N:�ɧT�K#e&h �t��Tƺ�8�IS3�RQ�	p��se�A5��+�j���b�-Y���԰:��LE���0�ʌGb�$ꢮ�K�U˚����(�k!1fW}l��q.z%H;~wC���vr�^�s���..�w��("r�d@R�
�@_A�	Q3
��!�c�ﾄ��J��F��H�O�A\���bB�b�L��>�Ppy������$]6cd(���U�;���v��$��0$�]Ph�`���� ���av��*�E#M���G$�+0y_Ua����Ւ�/_�x8CP�N� ֤�E��^jet%^�U��*	��
�4������(�T�Р�ݼ��Ech���g5 �bs@����p;NQ�����: pJ��H�Ӏ��ê(�΍��fP3��`AW��:T3������Ńh��axC(8�_"s {��c�!���s�Nx�ʜ  ��ȡI���Dy"�� ( ۾��8�>F��Ȁ9�UhZ�)ժ�m�Q��V��TZ��\�U[cI�R
,������Uh+�Q��TZ�M�E\�|��O�� -�<������������~��j.ݸWa�=l�g���>�����
?�o����������D?��� O���#~����Ѣc� B�s㮏1?�}�߈���qPä   J��R"- �E�v�bB� 
)QV�":`P �q�s"
�14���@*�R���w�p�D HH � �ƒ���E@�	 ��+
��U�X�nw���[7w�� �E(@��`*�PE�UJ�j �A���i! Uߑ\
 � dT� �����]�3�-5��Kw�yv�6�N�$�"RFe
�B{�M������G� �
�(UZ�]�cs��{�@��ә|,`fB���-�7#\i��ca�d�e�U�&,F���3bL�J�$��hg	�Q@�	fTh q(
:@�� JTDZ���(f̦!sb�lɍ+M�l�0d�N�����|0���R|2|u]o�4̰	�,���Zaե=H�Њ�-?�\�H������?3��uC�����gM��rw'{��$&,�Fw>�����2���|�f}Hh�ٿ�o[.g��P�ǟc	�z,\W�'{�K�
�X��K7�lT�&2a�X�<��{�}���O���,�;�ֺ��}���"��\�)	9����d���y��>ތ����w"�Lc=+T��{�R�Y��� /��(V)F[|*L�����3"���0���<5Ig��Kq�`��>��؁�J@����;��V}+$�%�$�M,�:� ���_,1/-ݦ�Wԓ�K ��^���Nbc�J%���}���,
Kg��f|D��<uaZ�C�(]nX�L�h��??W��>�!����c���cG�}e�H�|L�� �钑9O���b�#cDQO�]/��Q��䄵"U�"g}e,$cl�|���qKm�_x�R;��S�BmJ�o|� 1�>�M�8��K&��{Lm7Vu�$�3Z����2��YX	�����B!ORP�X/,����.}�	�%R��HG4&��?}���a?2±�ϏY�-�'�"�Z��g2�e�[��<L[����i����������#�2�ٝ�[dl�0���J D��ٛV�ܡ'���+'��θ4�=�w3<',㤵�� ���=�?��@�/ͫ`�)���<��T#z�J�� ��g���˵��Z�����B[^׷tN~f�3�i>�ڭ}jx's1.�Ly9�������>/r�/Їš�,a����l^}p�S�&T�(��5�d�j��O\�bS/���hz|��*f�V��3~���l[G�t��3�ʁ��]=���xj0us�Y���qe�Ա��n���V�����)8�?3����\,�k,���>#����L�c���Vu�biCǀ'̿/8�Ն42:YR�	��[�|�Bf�Z��m��}�
D+��$	5�ke<+[|�P.��pX|y$<�I�~(N����I ">c���qӾ��|ui�2$��H���MـaX�[�[}�׻������t%�a��q��7}�u=eS�MQ��3%��x���O�AR�2�!�d�3�>{绬�BT9h1�9e���F�6�R}��'�Z���eNl��ǌJI�ᵾ@��x&Y�U�O}���֜`!�X���-��yTf̟�>j��z�1������f�)'�5���2��n�������N=;!C����|0��r�@)F/�>�S0GW�޿��/�➜@���>��L����dTp��y����.��%c&�� �{�}��Y@'�Z�$�$a6ͦ��牵[|n�JE`(�	ǪI�
��;�� �!
��X1��C�b����̤ �HfufY�^bL����wD���,	�cJLQ&��%N��27���5��4֢{�����2���!�9���gW��(։(fk�v�)�[�]���*�g�qYvƁYkD1#�v��a���A>�R��to�f����)�깪F�\ �"��!��O�Ƿ�qZ_O�Bx!RD�'�)t�-B��?|���KǓ0��Rǈ�!>Z�-��I8�`Tf��k��*Ɏ�ۏL#Z)6�0�|c�1}o���n�"�P�X��^��5�M�Ca�N.#�wR�#�U�Z�Pm���y��s��*}��'ܙ�>���@����o���w�,a<�R�������ӪN�Hs��,O�O�,�;Ї[� �jE�P�U��7�ǩ2�l8��e��u�s�-���[�l����&\�g��)!���U��@�y̵��)���n�����o�8���~�Ƈ<z��©�9g�{�E�������N��$���岊%��/����7�#4��\�y��[j'��z`�i��a=� F��cOsc�b��ٚ[RZr�gZ,|{�h0�C���F����������^q�!�	�3e!_��E5
IVIO�ˆD�X���.e�|�P��X'�c,<>��gd�Z�X�C���)�[n>�U��S6}�K4��ӓ�#���XB��WJG��!��2���k6��;�����Ⓨv��������"j�r�H�u�'wi�ITA@����_�t�>-HqOg	D�'���n}�φ�~�}Hf�O�QB@9B=���Be��(ep��P�XK ��e�2�<{�g�ӹ�]ɥo.�
��k�O�p�&����%_ C,%t�_<ίk��Y�++���sau��V�� �K�>��,R���l��ͽ9��C�<G)����0���h��!�����ȯ�|!	 ��'�sݨ_uAnw�
�Y�I��=�%�|�>$"�dBfL�T�O�}���X|c��E�K�%<�M���HD@�<z��2}�����}P�3o3�|}�S��Q�<?���i>&���(B'�̏�6��0<��HPXB�<	O��4�Q"���a��N&��ZS���։J�I�g(LƏ8����Y�����U�<v��}o�c��|%�@H���|�n���)��� D|��4��$x��P\^ձ+��Wv���}�s�W-�n�����c1���R��k�H��{�*�\���ɷ6�.(R��!B�k�+Hθhs�&�榅(��|E�|G�x�b�b�Y�?�Q�$y�Pa�80�JH���;-�%y֯��Wzu[~�u(�@����jn�AD@i�w�3��~W�o�W�;��{�����ʇ��
��{��~_��<�'�J���*�I�
�����W�?�ُ���D�G8��������M�i+�`��#�ɯ�:U��6��4�=5��5�����k�J~P'�w��d�u.�����މ��{ݗ��C���#��[D�9�����l�X���5�aO=\#�a�1��G.o�����6Mc~1�Μ�&���j�[P�J�@@(�(��(bP
@QCf��1�C�x#RA:��5���b�nc	g�s��8��ݾ}��8d�.c�=�o8���b�~o�7��k��fc��4P/�U�$�duֈ�#D$����J	LB�X �%w�W,$�2�L D �!��A��#Yq��E���WK}z��o�`ۜ�[��^b�cI"\���w����Q�Fn��	��Ov��Ӝ�����bD"2+����@�����2�Ҏ�$����ݡo�D��s�2$�鹨ƍk��V�ͫm�U�+�ܭ�W�j{��ݮ/-r���۔�$��%�7wj�s� o�pys��"��%��wt���$����dnt$^]H�3E�#y\����I؏u�E^m�Dę}V��&G�Q}-���F��R���yk���梢�(��nr����xI��{�˖�\ƺy���b�ffX��Ģ4���3M����)e(�^{������c��f�I2 %�jR%*fA%$]4��+1���k��b��݊5]�\�ۑQG9c��X78y���_;�c>u�G:\HėwIe fwF�̊�'-�n��@��@�ō����I$�ܨ�sW9���|kk�l���z���.ǜ�r���wF]wH(�����4j1$Q\�]�ęc%IDBB0њ�шy�F��ί,���TX�5�#8D����{~����s�}^��t�����������_��a��C����I����C�����ɝ@��`����������6���o�Ϭ_�j��s�s����X�M?���%���A1f���#�A�{���Ї/�{�+������CU@�- �������d1%c���+����-��DQ�޽q6P�v�������M�˗>��ݺ���D)H��tI	���40��hf5����խ��cE#�&��k���kΝ]�p^:��-X[���G܍q�ʨ"��j���r�la;l� ��y���L4��P�XYr���
��jҮ�D��U{���OV�l�����;�
&���H��5�O~QT� Mo���)c"��Y�n���9�C��P|��i����@����V�o<�#r�DW.���D"�j�PE�$W.I���D.�HcLۻrn�r���ؒ����;��Rc`�s�;�+��`��HQ!Q��X��P%%9�4�:�@s*���-�͹#�b�u�;��g]�W7�I,(˛�w\6"ht��a��h%�H_A`ā�"��Ƃwk���{����1h�i"�(Mu�o���7��2������L�}�3�K�w�~Eqk_V��#
�`�2�"���\�腾��Rd<�A�l��NBpk�C�S��/����/�fM��K��je���$������)�i�g��ڋ���c��߀�Q&{��o�����@k�'��B"8V�׃� �
�zȞ��Ƶ+�4��@����{�I�ݦ�j	JR��&�$�z���uG{�c�� D�!��d�B�������Z��ן�8�	g�.��	�aᦑ��k�uL^nk܌����\i���L[)����LG'��ae�u|*�2q�^����h��+O�W�MK{�xw`��E��qȵ�ݳXwuz�l����}T�R�_�,E��t��X�g4(cT
K� Q&X�*��2��"��;*/S������]�m�5_����Ԙ*#U�e჊���'�8@��^*2R�S��A�����Sw�z��y��������ih�qKH@��hv�
8\�-����Rf�u�G��){&�lف�|���oS�W_b��D����������a�K�ѭ���y뷣1]���yvaW�%����W:��tu������~���u�C碽mA�����+�K&�7���F�!Qywa7:I�}A�����߼����d�b�/ͬC���ߦ����w�+V9������sߤ��N�댃H��p�.i%ȷ*h�;���u���M���>�|���S��U�rE������+1D��e$N�/[(�%��;����'^�F�k�P��H�3眷R������}`�Jᐩ�)^[M���*0���v=�j�ѧ�gs��5�y��|/�)�-�f"ezخ'r"鋥oD����4W=َ�R�>�a�nƽ��Q�L<J���D���9ʛ�!P��O��`j���4�z*��DgR`B��6ֵ����JQ\^|��-�~Đ�T�=���ޛ��^�o�9�H[�j��4�ʾH�2d�U��T5���+kl���ܖ�W��,#>Q3�,<��K*P������s�X�<��%'��>x�|��*M
���p����Ff��Պ{\���O�{�X_w�9�|;
ey��ԸV\���#u2��N��)K{�#��yQ�&����U)�Ȯ�\+�T��n�Vvԙ��E1���y��!�>h$ߍ�Ob��Bg�;w�%�n>����?�����1A�Fy�7��b8u�	B�������x�|Q��4/\�K'���$gS���a��.�wa#n�~lsXm�i|.���?U�R�B�\�����=��r��O]W���Q�Q��Sp�i}�-aP���M#��1�m7�/��`�Z-���˗�m��g���E+	K9�ol������6��N����S�m�>Ȉ�u)�V:Hd��3{]Zh�>���_&?]N�LXgQ���Z�*>+�����o�,Z~z�3�rw�ʕ}�C	s��i������+�&�h1,%iz4rkn�P������+�	499Rp��ϢT쳆9��Qx�җ��c�S(>�<�*�H���JA���e^�����#��Ed@���0�1�ɇ������p7��Ւ��<����مZ/U�������p��X��qgn�����QG�O�L��iZ�O��KDy��	�rh��u���ŖZԃ��ڃ�y��	����ƃy9����Wv�_*�o�Q�̖����w+^v�L|�H�f�o�կw��w^ƌڜ�M�+���/1{s��{��PR0&���Ѽ�d��㏎�Wz��k�N������T�?{q�_�]����\�3�Z8�1z���W�Xټ�������b�U�'�%R!��l��� �� ��d�*�k9���n����#	c�{�N�C���{-޼��U�1Տ�?��2�^��D��{f|��k��]�(|�\�O����lHi�t�b��Q�Cjx6D6��#1�'�޴U갮H�YDT*jRK�c�GP�ˉ��t���wyz��g��]ㇻx/�{�����$���1���5�F5��1�}��5��M�����X���ݗu;���a��3D��>9 �1L���7��u�gpt`���|�(�&0Qj4IIE湲V��[�ʸW6��-��5lV�����M�|�z��蘹sG;��ݦ^k���%�Jh;�f@̄
wU�wmԇ��.�du�43b*6{������,B�tcY7���皼Ѩ5�wj־kWmy�ۦ�4F�(�2!��9��u�@��U�%	)�/Y`C�%$RFQ�h���5�p�{�"�ؿ�Z娊�j�V�k^[m6�嶻�H�빻��� ŒH�$y�L��HPtA��&��bNvwt��]݇vƺ'|��	�\�/�e��T[24�E��n[|C@QE#M����Qr�z,�p��(IJ(�uw�IHH��&h��/+����PRY�U�+/v��ѷ��E�;�*���j�km�Z��+	��W�wt���	���Dw[�ʹ���c`��T�TT4RL�����q��{��_��D<����������������G��C��B���g�I��{���������g�I�HQXb+�/��;?��������K�`��$���|��`�c���s�S��4�C*���fG ef����66��&Y7tq�4��Zɒ	Htppȫp�B���뀕��?���{8����0/��$%`f�bͧt�U�����x!����i1L#�떏J�ui/��d�F�+*e��d&� E���M81�Q��R����d" S�U�ʇiy�5���[}�$�LF�@�i���ݠ�S-�E����A��A���z9����_u�PD��@�V�@ ��8Xc ��&�!E+�L"���?�|se�RE��4@�n'&!�VLxR۾���9>`�����	�ɠ�Y�+�u�F�ԣ�09�����UHՏ��/D���Y`I������h��/]!,�Iȡd�$A(6�(��SR"y�D�/o��p��!P,�00�@Ƀ���	��e`�W��W��Q�	X��a��vֹ�0!��` �(c�`m�m*)Y�&%��v�u��ܖA�h��KFF �Jͨ+�"���)�_�j�����8�n�c�G���:e&�Q:2.C�0��m] �$i��c�'�4��m�E�WZY~�(A�o�a�2����Y&r͛,�07~�<��Ȇ����4 ��l˱���� �(����W�۸�wf(�aF ���!F�����2��L1�m�W�C�4�Fp��F�t6C�e����f\�C��=ͰuϾ2h�c�Z�JX����2K��=2��1�qj���DH�Cڭ�,I��M�m���Q�ܡ{9�/��6�]$�:�2a*P�Y������� �_]3qP����\�p�$�e��T$p��o�x!��;�Vo����cf6���\z�5t`��\[J��;����ń>���>�H�'q���	���b-�&�i��&���2,ېtS�����(V
����<��t;11O���J�Ȩ����i�@���h덢H)�)��J|�/u*'�ǥ�4���G~�xPН�HjVMY|
vꨉ�,E<
����������+X�0M3ݕ�4��>3�\��jֽDH�5�hS㱤�����W5`�Ҥ�u�`�INi��%��d�L'����ÊG �\�+SBob�,��ױ�B&�ܳ�,B�P4]��S 2e��vE ���r��"ZM�CI�Ȗ�H�(�Ȩ�	fo|m�UP3�� R��ՠ0�dM�j�룐��
/y=R�b�J��P��B�F[1��<'y���ˁ�p�N�S���(�1��QK��4[%Ͷ���6-�j��֊����P�܄�w]�Ɋ�_�:& Owu�B�+���ذX�H�t4�y]݉��=�ұ��b�j湵Xڍ�I�y!<�=Y-b�������w@d�+�(��43�4���owub��h&Z��ƼMBm�]�#�����B8��u��'ǩ�&GκB�D�1���w(*K�廸)v��Q�cE��(�[�m��*Ƣ��r���FWv�F�����1%9��EΤAS�s�[��(�,P\�
"�$my���,Q�RV�ڹVƫ�����Cr�D�( h�s���%�/��&(|U�Q󺴒mQm�E���F�"g�M9vX��u`ܸE�wD�5����ubA|�QEh�j򭹭r�ROu�K�%F6>wd9vO{�j��r�����(�[�řE��#;#�5�ۚ,k"k&�\��מTb+E弭�E�ͮm��u�I���EI���Ch*Ɗ-�*�ko��6�D��"T-/V+�[%.!��1:�Ư�V�U}�\���tJ��sE�}}���^���mL�I|nXѬTk5�/-�mX��PU�_�^��m�9�9K�F5%t��ű&��F��C��Z�Zƪ6�-�+Q����kkn�}Ϻ��w�����ں�ޝ�wj�5�m�V6�\�nk�9��и�1Bc��������}s~��x��������������'�ǻ�����x=��~�������W�p�?��:�i�%s�m}^��/��s`�b�G_-
	U?E��Q�_t��y�P[�k��Ӗ��m�FƱ�"�6*�F�5�Mk�-;���H�������r�Z劢�}��msW(��fl[F�^mtڊ���"(�y��m&+��b�Q���u��k�[_�#F�jB�LQm�T[�-��b���sj(֍��EE�5sX��s��M��$����&�t�*1�km�[^�H!뚌�J�$�V1`��o/6�ѱ�[��k_���#F�W��Q-m&�E�WKb����)�Q��ĠR� �_icI7H#>u�k�ֹ�u�:m�owlF���ծm���m^X�kͶ�0���dń���4�cRF������hجcUk�{�3��w�Y^�Wwǻ��k�u׻����\1$Q�QZ5F�Q�j�k��[Q�b�򭼻���$%���؋!����ы*��
-��X���[��{�M:wE$�f櫧��"����)6��V}v�F�F#|nXت�-�sj�+�۷��w\�T��D�Jd�G.�����"�nj���1�r�Ed6���1�R��̀��k�E%:.l��#Es:�&"i�Қ65s��F��M�>���pZ65s\)hZR�����U� �3c�4[���U�(���r�wf �Q�F�EI3Q�kco�k�lj��5�R�����"��nW����9�6����E�t��I����5��s]5,j �2����ĉ�F�Z@G��sb�F��E��p����1�u�����'u�JR�Y]ܓI�sr=�F�Er������JAĢ���rK�4�d���ۗ��-�w"���Ԅ��N�s�wn����=��EL�-�M�6���\�Z�\ZA� b
DWT��0Z�5��r
��Fs�N�s�	ˁL��\��Uɋ�;��(�%"!"�6�m�m�Z��[v�o|�^TZ6��y˥ϝ����t�\�����RW����%��L ���\�A79���ԛ�V6�1�"��Q1"�P��QC
9��r��M�b��#nc��Ww\5%�H[wu�v�tL��(�hӺ任��d�$[˔%HWu�-cK�[F�⪋W-�9�C0
�9�B!bqb���j4�ʒ�uۥs�	4�IIΓ,�s����46�ŃD[��Q!�E�t�D1��3)�O���{�����Oc�g���DM��5X�cguvf$3�a���f�s��2I4��]��H�ܑt�M`��"���6�ؼ��Uʋ���-F/��o�ۦ1%�t����l��;�zG�Ǚ)nn�)ݺ34yv�	
5���m�mQi�8�(P� %
��\����j卷-�-rE]�k����/|�!�y\�r^\#9�i9�	�:�.k��>N��sC���Q�H�0���|�F�L�[�{�b�"����4�J ֪墳�Ah�
�������7L�"2%�sk�d��f%! ����#wu%�Ɛ�9�HM�tEˆS6�����mm���5�(���P��P�L�,TX�WH���ȭ�\�k�E�ʍ��ʦ|[�	y�Vg�ܽ�jn�5��,I$.]J����w0¹��va�	F����Ɋdo��[�k���͹��w�GW @'�R*d��H�6�Dh��/����l��O��;�g�޲�=G���������=������
(����W�7��u9�͚��E�e�" ?�{ϴ�O��_�To�{����W���^�������?��D�����{����?�-���?���e����MYO��_���iG�]����֤�?�N7��7��LI_��C����a�o��P�?��Y��z??n�   �5[O	�DH����g�9��o��"�L�B���W�Sr�Ϛv��r�˽e" U��'���=��{|D52K�ߗ[�P��?S��S��h�z�F���.���?�gDo������k1��i	Czǲ�r"�VH��Y\R�A��}>��4�	�X/�o�ri��핪\3��$��K'�&�z2NZq���Y���&�a�}�Єd�W���BUY����O��)Y�c7��yOª�<?��iwBn	���Z��%�'�Q�ڣd��JF{��V���[3��U^&f�	�y�P�;��ںsW���u�f.q+am����bS/-$2�P����U�kߎ2������m13�|���Ϗ5����][�r��|m�;%�])C��#��:㓦
yMs���2T��M�].�,}`����x(�ŏ����a���Լ�(�Mf��p�ڞ��s��5�6����7N��ۆ]�R����`�>E�,f耸��HYZ��X�b�J��̘W(QAr16�3�J-�o\������=����r�"�б����VTD�xK����4Tv�8y�x�T��'R��&E�5!����رL4�B���[|J
��!��+�Ն����( "��oW�X��U�G�X��� ]�X$<x7�8d��������ve��yu�y���I_f��X]+�о3����+�C�I�.��q�2�z���H�6���_�I	U�;'�p���y�*k���rhڈ�v@b�)M�Ī�E���c�D�v@W A��,�ӼG���{��y��(�-w�j�������7=M��+U���I���b��|C:.�7��DE��.��̈́u(CFׅ��ozv˩�h��K��:��B�V�k�ڽC�GYW�(��Ƃ�w7�S��������?��[-���X3?�]�x�2Sd�]b
�;�_k:�snNd�)-�L W��m�-/ʾ�:�u��'N�-����nc�y��2j��q �v�ߥTn�BΕz�D�DJ��2�Q�����'�x�+�Gb��D3�v��y�}�j�Pr��H!�(��
�m���^h�{�FT�ߟ-]���Ѯ�qP�p������ ԅ�)���yo�k�Sk�w����Qq�0�x�
*,S��J��4C84�/#���^�i>JY��"t?7��GXyR��-���Kq�sf�k|~^H{��*�e�a���WX�KUw�8�馢�8���X������d{�_ �Tf됮6����/o4?�}����)5��Xg��&=C�+�����q3z�t�+]5B�v͘=B:�Q�s#�On�Fxdӝb�f?=��C����Znؑ��R�#�g�Gȱ���+2���$����K>���.T�1K�t�4����
Ct���e/�Hkg�{�$R�ACq{�1�7Pq*l����N6�V��m˫廬=LY*����|o++��3�i�~��/�i�h	M��>o�!�kO,���:.�+��&t�[$(��6*�R'�����f��W���j8�`TT�K�:�r�h��C�Q��+W�}aHfb��3�2��Mz��E���u{ҍ �m:��3���5'�:�gƦz�Z�@Y�U&�vjWp-�¤Ȱ�RxA=0��ؑ�m�S���5@*�1�#������L�ND��6h�y_k2�{o2Rn#��� гq"?6ƞ��x[�s/�*F��@wH�墠E@��`��ެKE!]����A���r��cی9�=��|	�M4���nz�*N`^SIk��D��e�c����/�#n�Q��}u-mnw�k�nӘ�]�T��k»w�f����%���OÂ=��H�����ɼc���m� ����.���Q[��+I�F���g���_��Q!�����w����ӕ�G�h���I�vQ����,j���8�6T���\�1X[x�����ۋ�%w��N? e���EF?%�B%���jf^!�^��i������&ڪ��~4V1���#��%L�R<���X�S���:�~XC��`�k4|@�M����'"�WJx��N���
AJ�q��m�|9u�!����8����߲��x���H��ز@��M��:=ƻ�7c����� z��}���������}w���6�����[�}��n'%^��uo�7vJ׮�m��D۷������w�;�[�Il���#.#���L z��-��e�$���H�� \���$/�������"�%�����Nt�q��������Q��+M/�[��.�l�Ue���?��0��X����)R��	_�?�,����1�O�R����8E�AJ���uci�?�M�o%#�W-�[$t���OD��Z"����x�u8�)�aE3�t����405��fff+�a��t-�9eU���7�5����fB�<ͭ��� P��A��`ؤ�WQk�@u���@�E�Z�/�3�x,�4
[�ͤU
2=��Q6�J��ڲ�>b��d>��G��k]����Z�N �dDCCIh��,���Pd���jhW�#Q�6��Z�ľ:�c�-�) �����݆�rc℉sfq�%O�hG$@º��	p��'Z����W1�y0pE�twy��ZCI��5<�;M6��^��
Xo��y������#�QQ6|�N;�4p�y�I�EF�G�	�%�E\n�4Tu���LE��R�	E�x�&��B�(a�d���(���@p�$ps�BK�A{0HdE,@d��QU�]��X���5�+�m�HM�(Ac�p��ȭG9v�E'�q ��N<��0�N=�L����}EU,�%*��|��IM�A���&�o� T�hj2��>P����<B������;�V����شB�(�K"`F� �9��2n6
RZK���n�2,J��QA��#�07J�%��[q�,��	#p�ʉ�Hw="A1ɢ�C�Y�`�%A�@�ϔqS@m�3���P���ق"≔c�b1�
2K�l�%@�CX��E#o7�V�r��,��k1��U8����kOx���2bT�[95�E=��4X!��v{˲��,��L�ӯ��]=��Xғi� ��
h�e;�VJ�ܫ΄q�4yR�p��y�R���\R��T���KS��<[�U��x�NV����q�c����+ �q*��ھ�f؅�2�@Ue��ȍ�:͐�1B��W�7l�Us��96@ۦ�r�q���Eh\����~���L�\��q��U�I��������I/'<۸X5����d��؞>M) �"2(���i����b�:d[�:$"P7!D�6aY�6u�7�VB1D�H�|�n�w�j�s��|�.`Z�  1 ���~`znڐ��`1biV��J�F� �Żjm/7ko�����^;���M�x�C菢47|v̙�1��j&�6fP"�*mlV�-jJ�҈��x@L��h ���� @���������;�|���!��9�@O�1�?�}��H�S�Ŀ0߮�������de?���������������C����_�^	�%��O�E?�H��Ai�;
'�t����%��j/続���_O��P�y �r�'�ɞ��b����J\��vȳ��izO��O�w��O_<���:��Sn�����{��m�P6�E6��J��o��#���I��.���D���w1y�?3BZ쪌�1yL�����\OqW=�P���oH�^����}уk^ֽ�Nb|� ��>�@������V�7�:2&D�2a̚F|�6yGO�*K�\���<��P����%��f��D�����Y�G��\j�|Biٰxk���,~����>�,��և�(o'�t���t!�㠑���S�H
O-R9�)-m��
[�F�y���|��~��t΢��������`��Q���un�����%����`M��ܛ.��,�;��H�������v;�����3�q��C��!,��m�E��eB&@�o@Hf�qc���`m�3�i�^�b�����Q�o���l�j\��tSs͝��-��!nn��f7�`uY�N
�m굫��e����EY#�%���X�ח��tf���	ۀ�>q����<(��X̉���c�Ķ��=�aŗ
$Q��^J���yð���<�-JS�i����m��;��w��y����Vy�(�U]#�L�|7�L2h�'�؜z�[�l�Xd�~G<o�_D@��Q1��g�Bn��6��VKB�3s,[}t�� ����vT��� ,��-��8L��1������&^��0�>�`���mߞ�����D۟8Uf.�Ì���lF{�q�{��ID��Hd�*2l���M�ė�nxE�D�3��zX)��f�ٱ��?D(�t�є���8��湆}��׸x4���L�H�_&K4B,6����z��7�aKz���x�s����3�*y�AHa�hz>���"��Y��l�rY.��y�f��Ba�r�E�G�5��W�̅v��ov&������K!�O04�,�E6�<iS��K��x�Rt����ؙ��E-t���[�M}���Ԑm��@�^a��>.�籄��b�^:��'�l;6�}^rp^S����a�)hje����i�'v-c���+))>�qx�K�{����Ċ��^��^s}��3���Z�T�!.��?u"��m����=�܆m����"�h����e�b�D�����W�]/�w��+}(hy�*�}���V=��38ڤl7-��q�B��wNq���&�8>���<pV�c���J>��E( �|�Y,�rXy�tק']	��6��N�^������h�k7�70�`�b��z�Ȼ�7����Uw��A'�0'B�c��\�UXzR2�J�>�8�5�W�����V2��.d�t-��7�h�t'@�KI$��Lq/����^��#��Ϸq���&�C��h�:V�n�a������^z��H�K�S���󝫱;�6UkkCo��&��D� ��w� ��y�\�K���朎�����u!�Xy+�1���r�jA�e�_R����w�ޔcR+�aգџ9���ٽZ�FO8+�NӄG}��J7��ie��Y"�y���+lJ�~c๛�j�r���^ë���'d'�KR|��]vw���G]���g�م7e|�D#'����q��qy���m�%�Yvde ��#����F� �
�`G?#������*�}����O��6^0D�r�B�-�c['�z�|5%��\���Qo4����D�ˢZ�;�DG'M�W��(��ǋ���[��E�4OM�7`vƶ�گD�zj�{�q�\�_(=�{�d�u�;5�q'�8~�ܕnW\Њ�Q�i|��k�NG"��-n�p����$jz�69���#?<�I�$U��{>x�0{g���cg�1��x��잧�v#�hBޚ�+{K�$m{@tZ��7����r�3�ċ 3�;���B��s��a Mb!o�[�R�܆ l@��2�C-���+=��E;�s��<�3[�V�[[x��cuI����/S%�6��|Ȗ1W�X{;�j���.�.��7��O���n�{�<�z��p𢘮�%�Ӕ��I�Ihɖe�׳a�qQ����~�Z�5����x��FC\�'��?N�K�-�T�K��/�v���O�>�W����?H@@� !�����_a��k�k�F �j����iբ������[?�1J�G:�n�y�����]����5)n8�~����~*_����T���j���?u�h���~��$(���q�ȯ���<Xg�I�=C��$?��s�o���r/"H�3� ,WUQA���W�8� W�RP�ܺ֋ ���`\@(�����DT���9�����$AP`�N���ơd�i'���( �#օ�x� K0��7h��'}���� �L!5���kV�[�PeU�f�#
�Z�Z�2��5�:��h�0�$Rxl� ?�d��"7Du���p�(T(T"+�R
��F�zo�i���1ޙΞ�Y���Fe邃�t�KȄ��1P��݀�<B�,9]:�M��jA��jWa	�x��PW5��f��l��.sS-�F����j)�j�x��鉔&�B�"��6A$us)�+xJ�����J�ĉV=t���O������h��^+�W���;,�z@��:dZ&�FF��$j���|H!@0S 
�R��'�S&���*p�̰�<r�!]уAoP.BV>! rJ8�PԹ�$dB�e�N:&��X��%e�
�Mr�!Kȼv
D��O=���	
� �����EGl0���i�m�����S��]!�Aa�
Ҩ�"V��8��q.d��If6ь��˼\�&]G)1֔�+�m�0�`�8 B���Ld^���al�j�v��yZ4шQ����DH�IN
��E*-�,dG{B�u�Q�S
@�BdK08�@'�Ѭ:S)z����T�I &C��0S�,	1�!�A�(.�mW����-�E?,[|.f�F@�#%������es$�ȩ�U�^����]#�g/UޤADx��]�%��%�����6Q9�k��jo��䗛os���#|=&�y_�p�x��̑2�r�2Cf��n澂"a��i���$�DS���0���/9,�f\�+����gYlϐ��yM;�#����������.�		�j"$wچ�0���<�*,�P3���\���`���DA���'!��'t� 2�N����6��H�3YZ�ˍtd��K���4�0����U�7�K��&rn����y��/o�_�@e`�?� Q�2 A�pQT�Lض+]�@�MF�4ͩ%)�"d(̆�(�!�_��o���)�����^0_Jx��<�DA�F`P �Q\(	�@T! %	?�����_��.?�����_���'��G��W����@����c;�f4{���߻�O�D���~%��D��(v��������ƀk�EcG�J�˫���C�_���?	*誣��DE���4�a��k���I,��=au-������6�O �N� >��} ���nO�������E�Ϟ���3v�˙X
� ���~�z����ȚV�A�'��8g�Fkx��,�Esҙ����t��`�y*�hl��;��+/����۽�}Y��ڎ�"�S�P�3�l£h[i�۝�=��R��)%$$��t�����~.����x�Q�j��B���W�w�n������� q�D��=[�y[ߙҖ�}�g�d���~��8��.꺱-S|��.<�n�^�=���N*`�
r��<4����O���1"y7vtV2`��aE�%��{�7,��*r��\}���Yf.�����~���
?�+�~�KGcN�����5y �����ԉ�]�3"#9��<�vU(� y��^4iV��箬�h<gBȿ�u��*��yڻ�n�	�F�!W�V�<�7kǔ7���T�ΐ���/�h�<�nm���"S�^{�+�LٗlN��Z�(v1G<d�R{"�.�ޔ�X'��V}"
�`}o�)f�ڇ��.3Gr9�DiZ�N8�;������۹�i���1��Ϲ? r�KF\5�V��d���W���t�РT*#W��&9<��5/�:�p�vH5V�b��~G*9t�+l�}R&Y:G�Ee��!ɑI	\�m.)-�{�&R^�m]ґ�w��썚�T�E.�f߲$���q�okFVJ�O��:*GB�D����hR3�}*���q��~)�+8�sW�rO����I�nm�b~Q�@�@u���J�ylb$�c�{�QS
�|5n��Ъ�>E=�3�jq���&��(��Qk����A��X��g4ǋa<vs������e���%��o�0F��#�Ǿj��S�]^ɡ�U%m-��ыx�8���/[ٽ��������L��{�0�Mw5��8O�z��u8��a�o�R6�ZN�S�щ;*ut5Y�n����)���1۳/�U���jW#<8�S����%���$�v�7��'�ߤ]�� ҹ�o�X�3!u�ds��*�3��t����W�_S�)�W���-p�9���$���lЩ�2�L�Y�Š�7ig%`�=k�\���_&��3�X���R���==7YwSW��P�a�sIx�mxۖ��w��i�L�O5ZB|]�3��k�C�r=6i�j�;��ɟP�Sl����;��^��{J�C3o���ݭl��i�.]*�㫼��:@ӫ��C^�?3��ի��`�}Q��P^���Py;�^�>B��n����T�e��������Wa;�q�c�{��ܯ��J*21�i�f�|q��7x��[R���?�[┴LweeO��{��,����7�����v��\��G
�Œ������k�=�V�k�иt��8�%s$z��(��5�Yom�;���2�\� TК�6���������K�2D�r��FSN!l�)d
���:�AM��F/���h2o�$���H�$S�2�O��jC��v�4`�k�G=��|)l{a���W�:��U�$���9��P��+c�B�0f�N#�x�ة�a���Ng�'�O��/�v�B��m����_X��U��x�/!Om}�nVOy�T�h2��5��Z�\�-��e55��N�]8�����F���p���;H"ޜ#��hz�
40�R�.N��঴��E�沩�
g�VG(�Q
4c����Y ����`M��+�]ͨ����3�u#�O��B��tޙ���ٸ>|�[����V�Pb��-HHd���$���R�N�/&�ϊF]�}{�C�t�Eӏ��5������c*�Ze�an����\b<��F�������|w>�:0Ib���"�־I�-�=�uj(5�<!��U����@g�3j�K�7/x���_A�?&�U�qF�j�խ�1��d��f-�w{7(˛��󪿘y�NY�?)�f�����Ӎ?u���/���L����f)�[���� ��8�����#`��2�������DJo�"�ОD��n�-g�v��q.���b��\��'m���&=���X���		E+b��	��g����w���v='miฎ˟�pqu����XB`Y�e�{�����)��<o��/��������>q���*ݯ�����É�Tɷ������?��������$tߣ��F�з?�?V�2i��x�V{������>���L�~��W��;���mxQ6����p�,�Y|e���Q��j#+lо/�Z� �m�m���i�Z8�����i��S��	 e��U+uS��I��V�i��(6�-�[�>�e�
X���M�&��jR�TAAH @�ye�@뢓�\}4�<��y�-a�4s|��IT�-bG#B/mj���Uj�Mqp��������Ui$Ir��C.��_J��4u�� a( l�H�� ���%�zM�
H�`%㗲����7Б��P���$"��sTyBFC/��Fyh��q$	D�Zf�%1\�I2�ȶ��"U�MEҫ�MrM�F%h�^b�>�u����o�u�9�
6�I�g߼٢ZѭV���L�H� ��*��~Q�)��m9�6�D*[Kŏ|�,��B��8V=UM2�m,��M;�
�O}SN5�B@�$a�(�Gb"�T`0�ʪz%	D����8�p�^����H{	![Ʉ
 ��.9��F.�j��G����a�I+�}#�ڬ!h�A��$�H1B��&�u�Z�`\��&� ���A�=BF4�8��X�Q��1��"��Հ���D]�@a����0�)h�閎ID�Y	A�)<0���FE�t�qC�Q� 0^q��j	Q��54_�?�Mߧ��ʝ����s��ԑ� �������~�m �AU��	�� �oh.Z�p�2��B��)w9uͷA&�>	>A��X!&DP�@ ƨ=�E�m6�!AAt2���?Sk#L�+p	1���m��,>�$8�[���Bh2I�
��#-L�Z�kW\)��h�GXC�!�f��(�����w����(IEiVM
g-�<pb/���h�;l
�A�P��1S�I�Phힲ�b�@J�6�I�I�ukB	OY�����G�A�Ky�<�uZ���b��ڰ�Ȃ�E	M�oT�p@��w���n�zm�nϑ�gwߞ�,�JU�I��+���Z����ں�̦�?��?�Q_��㣾�{�`D���>���{�Ax~�}%��s����o�~�������~���P��M!'�����������?��%B�_���"o������/����ٸ'�o̔)��{�Y�ŝ��b��?�\l�]�u�	75uD���Jv���u��[T�;dޢ�RQ�t�ݰ���-���-W½��L!���(v�J�,��7Gگc����eJ���{��!~}
�lZZ �d�j���Ü$����f@��"K�j?���u�e%0oIx|Tw�%2@}"�Q�<���\������~~wjJ.��&�t�_w�� ��o�x��V:�.,FTj�p�i��ω����|��̞�C��B����2(P/�ݘ�-*�R^�T���MX�V�ҵ&�����m������ϒ�y�;~��!�؛=������t&I���,��V�+M����N��$�Pߕ��NF��l�]�G礠ڦ{KT�0�ަ���xJ�����^(��2���J��fs��势S8`�%X���|V���yG-#5X
+J�Yl���k��m��i+H�4�@S�%���ܷ�}�Z ukl�%�����j�в5�?�rV�*{�K�>LU~2��s"X�T�]�6����Uzg��)�%}aKy���96'��4��,��d�ك���c��4k6	L>5����e�M�:��y�o�x^9�K%�����!Ip>�=��L��h��\(��[�<��!�%�y?��05�yM+ ����m!Y��c�<��!���du�B8��E�#�4>`}jpk�ZЬ�V ��v/C��uZ��~;M��ݓj��VG]~_�"#��]I/���\Ѐ��������\�9�|W�{�-��MT������}.V/�ԏ����Ûߺ��Hm�V��K;�^%}"��JIAѬ\����e"S�Ĩ}5ۿÒωg�ৗ<*�To�}�O� �"���>�6I8�ƅ��=�9��5l�Ӭ��VcE���hx%5��PGν:8�k]����w���á��C�4�z��^co�*�O�v+b��ww�d+/D�FXK`|tr)7?��6f�K�yaB$jBI���ފ������Hل��yu����r��\�X�ء�Hz&ݷ�lA��w�I�u��[4�O�Y[Ƕo��H A�����<���{jj�F闍3,�	i���V�!�_;����lЪ�����R�{�Y
�9�4�� �j�w��uf��=��	���0C�h���Y��!/l��B�Уq�@_Qa�Sæ��L�{a����&�j���׵G����8�6�>�q4�*h#�g�~7����/��|�g�=���s��~�}K|t�x���^죲�R�^�lP׳���%����]J�ʲQ�����t�@u&�ј!�e�\��G"�)��	���߽/�8��g����G�2mV8���.��Vϻ���F����YE�ŝ�|ؼ��������ۛ�5��jYE?Ř]B�X��P�V���bgw*q����fE�R�6��$����My�'��bz���8�m��Te��h��]�>��eH�|�������]�DA��U��']gz;q��#�Gs�������m^�]���G�]����6 ̎F`E�U�{�7+�1I��n��Q3��9�@:�E2���G�K�����P�g(�	6w�⺶�}~����.�*`z�Ȥt�R\/�1b��lGbyW\uK��_��Ju��EA�2�z���ղ���U0W9�R�8ȶ��b�5�R�0�>��p�+y���5Zn�0L�V����7��省0��d�o�Gp�/j��˞�-9,|!?V����(S��μ�U�g�D>�С=H_�u�ᰖ]�?�4[9�fh�A�T�EY�w\d�-t훢�6���@����Emr���֔��Q�%z���d;ٺ��{kk�^ˮI~|Nwr����R��A�c�־�8���9��/��T�#[&_=��L���7��󧳿N��1�"��i�{����Q�$d'f5)L�.�4�v��(Ɉpy�_V?,�v銴�<%�ђU�~�!,I�k$�w��|p��Lmjg|�<=�񻬻��U��u~i9J����ۮ�Ce�?Ecee ��w*��^�'�$㮑�@O�׈KbӚD%8Dd7����r�p��hy'�}	�My�񲙒�&�D���@-������ͳ�v	%1�k��3�׮�a΢u�H�2ȏ��з�m�eo�OH�t+uiܯS���h��F�ѫ?H�u�>�}>�@}>��~����e}���߇��Do��?lS�;��'�+��O����s�'��Z���1U�@���_��?qr\���(T@�nH(�IL���G��<e/n���?=��cC��i��|�߯JǊ���WX��	R%C�C�	"@�(���)�A�(�N��L�ÆD�0��Xp�a�U�ʙT���l�E���*aI��*��!$�)�H�)Z�:�H<�I�Z
Ye�D*#6B �ڤ0�U(���� ��%����A��x�e#�T�P,X��B�	e,�Ә�O֪��XB�*�F"�ԙ$�Ѓ�p�@� ��Pah�0�X�«���(IR�&?T��ACPh�"Y-�� ��;��	J�%Z�����J�(A��a���Q��˒*�#�X�������H���ЬCQ=�g�(�-1��;&	@h��D�M��
(�̨��T��~�q4�9�㢭�ARDtҒ1�x���I|�p�������bd�D�if�%�JK�Z��y�00+`T�N��FdhaB�����	��-!(��	�T	Ѥs(�a�|�j;��ں�viw�Ο�9؝�Gދx���p5tj3N?i���%������;�>Vi/���Lk;{y���v.��5��²*�P+��vjG&R��G;�rm&:o�d0sD��H�5�͊�!�1b˼�QЙh�,�@ :ǔ�	��m�6�u\|�_z ��~�{���߫�q�Mw�ڥ�����`H�P	�R1�)#�*'�9ߩR�zrZ����(I�� ]��@m��lꝥ5���h%&�!$�Blg��Ի�,P���uVA�bc���p�_l
����i��'��d�[d�J��`�)9��El�cM��L��1'���*� b�Xt)&=.DP����*�)�Wi3	�eD�B��5W☙g���o]�t�[�F�I�l����V�ođ\ER��]��*��N�\�2��6Ҿ�Y�l$h�"i1�^[�z����_�_EĈk���q��:w��=������2v$tS�/5v(��3/��xs�j�jJX�S{�̫��A�5���͛;)���ت*�6�wd�
�0�F36+S�鼾��)`C]����KrkCº�v�R�r��l���<��;V�/of.kiI�5��˕�o�e'3��E2��'��pk�WgL���2%a�-�龹�DYp+%���[����jk�,.������SQ�*��e��t'\��[�3�Y��8��nl�J+�l&�¦�.��(U�L����^����h�u���d'�[�Y�S��E�ꀡ����E�0�����Ƚ�>�.Y���WS�l	���pF��Q�2��櫱˕�ջV��+��7ѸH.;��|�MC ���N���k'�⁁s�:���/�MV�s]�<"��|'wf~ϬX����Hl�H���L�lo�:^�cv'pD�X��>��Ꮂ�K&�W[���/bn�ls�Q�V`�V+~��e��:�d6�+�7�����r�:��k�^����ݑRrv9����s��)���s��輩�y��VNb�n��α���T��Sr�����B���T1ۚ{���[�e�0кz��l�����?�M��VD��x⹾��5�^g�y����o�/��D��&�����K���~��k�7�K�}u�@��'���)�sf���C�b2~����E��0z�M��4�������Qc.+��P�ߺg߯�K��!�C�	�}��\��#�ꤙI+R����AoΦ��{�L5��M#�<V��n3�=٣��"$/�oǷ��@���#��_}F!�ʉ�ў���g���ӥ����w����vwd����\%�u�KBi#N���ۼx��?�]�'	B�����t7f��}>�O�b_��rXه 2嶦yJFk�C�aJߌI���vl�#{W^={�	����3�Ԗ��]nz��P���N�Y.�8+�B���0�7�5�,q��2��q����mِ~���˲��R3�j�3o����Å�jo�X��ǧ����A�B�Lm����=3(��4�Л���d�w!��"�� W�]m��P�A2r%��5N��Y5�����@���%�cT+$�|ݸ����8J*����KѾ���\�.3e���7F%�	�±���fE�Bʁ��A]���p�YEÁ�_i�z�/�(���N9b��@�ӹ�Kq�X�R�z��"��^iP����%ua�i!�IG)q~0U��#=g�o|��_xEP;�[�v���osh���5:�����y=��p��g:��D�r�n�-qba~�9z|B
R�r{qL1���Y����5[�s&�%�;�S�Ne���U���SIC���>6�R�\�ae*d4���G���"��gt�(�<�Z/�����²���g]��{r���="�;=7r�K̎R���-*"L.���l��p?df�h�	~�Y���;�J%^��c��%�K�mz��������ݽW�����;��,�d�o׊l3�S�qxԑ�<�hP����JP\�>�~g�WH�Z��&|0�O�iE�@͛9bPp�M�/�U�r�N]���!G��A_�r��H�6��~{)���!��H����}ʋ�E��z,������ni�׶"��;0����2�13���Ci������"H�a�f�sݟR��*^����jV jjݩ��6]�rD�Z�����uЁ�s��~����t�j%���v�nLDȎ1��uj��~8͍���Q_[�+=<�3A�Ĺ���$=���l.>����vVE��t_)�d[�a�5�)&9���H�BH+b����T��m�*(��UK4��=y��� ���g�&Z���&?bzZ,s��*��J(@G|�V�2�����ę�+�Ƨ��}K���`�Ӛ�0]�iE쬞�v����S���)#�4=��P�������Ź�6}�O1�$iƆj%]9�}�5�W_�Z٠� �
��|� Լ['Fw/Xʳ3s��dG>�Σf�{l�n��l�e?�^�,���}Dd�:�:u���vv��j��^�'�6�L����>�6%��*���eQ��.��c1���k0}����#��w��V4l5�zK�E�ܵ���X���n�9]��_��|n�>
�rQ5R��ήQ���j��?˟�p����42v�\��vS@�Zcm��wltV�_���i�<��$��m�+1�!��H���M\�n����\����<��趺�m�/�s���K2k9Ʀ�VZi�����qbx(�B����������	't�e��t_��A4��:	Y)��!�l��$�ĸ�>I}wx���O�RA4!e���؞.j�y���'��z���N�U�����2׆{o���Q���W`T^�C��|iT~�ؠ�]vJ7�U8�a�����*�t��,��*R���=�A��Ү���~�c���NI*�iR�+�a��@���3]�'����x�$k�Ec<5�h9Չ-�5�|$�=�A<��QU%��h�}@�u���**_Q�W�bɋ�z��(-�I��{*7�~uA�!�H�\2�<4��Q�Z�?k����`S�㹯�;��͛T�������w�克����GW	���gK��j��[�'ɧ_2�;�ف��W�S�.h�;���/5��g�g�5�'��VN����a���ph�=p=�8�Yz��[mg�ERi	������"�8YggJ)��=b0�]�+��=���Z8c]�pU�"R�}��va�~���1�;��k�\���]y�$~�#�]���ѧ���ӻi�t��*Ė���"~B7�W[*��8�UGt�LOd�<��/�:h0{��i����_@}>�O��{�	����a�'��l���_�O�� �P~�'��i�EU�R��T�A_�P@_�1!�4�Z��pW�Օ��������-kF�g��^Wo�땙����r��8���C�:v���:����x�'�����;Y�Ͻ�?�e��fq�G~���S�xT�H��>'MǒK���-�4�9C�dT ������$�a�*���/����`�4�n�e1!��%�Ǎ�QE�����;i���ҵ3q��2w��ܯ�f���~�Aړ�qO�s�)-0i�0N{�N�f&ژj1�I,�N�M`"e!HD���gpBc��n�P	���gd��!�LiB�;D3m�2q�2@vR&f��Y�U0��t�ׁ��(�	I���5G�����<�#����w�4E�w�<���ʙzB5>e�'@{00�Mbc����#�HYU��A��R`�CΫ�	ډ?��ޢ3���7�m�-ӏх����������e��z4���%��(��!4(qL��8s�HUB��:�J@K�c@Uc���%a��*	 J
,Q��1���ǫ%����Vo���wjR���T����ʱڪ/묌�j
n��a(��~�}����{~����y$u6���R���ӌ� ��U�.DR\d]���
)ff$rɔ��CQ:ɠ'��7x����r�����ů�����#�����kΞ�Z	ac�-BK:0����zĮ�-L�G(䜔�vw�\:�&Tӫ8�J ��1'��Hu���@H�%��`���9((��B�$\�@	�e��>�<��bX�Q��� ���XL@�P�*��a*"3BB!L�I@P�;S��j*��LXX�_��������ôw_�׷�����[��|�w�$P���_[*���F�%���Ē�=tPj��_{��*���������Ӑ� x�[�1�V+ǟ���NLӟD=��Nbx[�Ě*��w�f�GQ9Q��i�MFڨE��
��[Vky�Z���Gt�0��qS�/bH�B�l��jhE��%����{ß:ڝ�ML�ѳaPq�i/,V�� ]U6���\�3$�.�K�aT0�g-�k)[ެ7M%|�!�[:�e\JV����Nv5njˎ˜�Im�7{g���ɍ9:�^8��H�c>��	�ø:F��̽�M�QN۷TVI�=�N��G�:O����Z��q�����fV�@Q7L���W�2���;6������OXrz�/6L�.���x1u�ʸ.f������mv@i���U�j��F�Sꓢg��o��T�@0"Yy�p�:��Mdi �=��w�Rw<e�f+��Lv}��\a�\4z��
c9k?m����+�9q��Yբ�Hv�TV.�ꍺ��Ȩ���Gnݻ�9r;�HLQ���'�W^XJ���þ�w��q�l������..�KHev��1W�^t܆v�c)�L)�&�E�qr�粄ew��h��1^�#� ���^{*�A�Վs�}m��[��q��p*//c��U�]ք� �Yl�=�r�� ��e���B̾��g�5�t��G@�&�^X�w!j��^�S5\���DU�˻�Q��m��'��#����	D��]J�n&��L,8el�t��P���w��> ;=�i;�\�¹<�t��<.���ǎ�����5釽���^�FQ�U��/̆#���\�[\ޘ�$^��v!�:3�o��e�k�L�Z�S�콁#5]���+�hJ��)�(�l�Q�]=�*r/ �ͽ�i7Z6_�qw�]漽�E�a�w�ﺵqY����۫�����\\�m�!��"{x��U`JT�\�9�9���_p�:!�R8]gL妮�q�t�ۻ�n��D����t�>o���/9�;�y�1�_9�z������\����������C���5���������?�?��&�+�}����zJ''���C�Pg�����_ܣ���~ǣy�c��Yk�������W��d<UQ��� �i����>0��.���B�G��j[��H��O�N�#�т��?q�u�&ɸ��=szC��$GCN�?�T�����!Ȭ���`�VR�uc
B
HT5
:�o�-$|y=9�Ј
���V[����H�c:%��(#J�Z'����?� O���T;D��8�Q����j;���U�}�h��$q�7���<��J���SWܿ
���?���ބW§N'ٗ�
BU��B�k|�Է����$SD�)�6	�]؎	�%h*-Q#��f�j�i��uIOJQ-�Y�
���dzfs}E���P6��j�e���}Hw�I;�]�Kk)b"�{��]G�l�%Wճ:��!��5?H2N��p��!�xg�YgB�M;����#ٹb�w���iHS�d�;��Dv^$Q.���qL��y<	��k��=ʒ%:7?�v�o0=�u�%���Ԇ]6�_��	�E;+H;[��6�'I$�c�\��1�ӊ>��N�$�/�i��h�{�N�Yyed�N9��ZKH��!qZ�cb�:�JW$aή�n��a:�A<���э*xQP�ݎգ��+1b��~A�nrTJ&�V��E6��.W�Q��#\'�쒪��D����
\���c	�;%��(��A�c;�;�Z�4|��]N�o�Gb��|�S��H2wwI����=S{�)[۹����V2Kܕ��3�����=xV^:1�D����z���u�����f��8}p]��Q1E��W�wcQ%��$�G�ݟ�W��n{»���}�^d����&!b]a3/��M�Z�.�&;���P���5{�u�	�̔',��b���\�Q�Nǿ�-���2�<�D��B��bs��x>f�s�wZV���A�n���^V_xE���Ps��|LҔȠ�-:C�
�M�m�d�b�/���1L>�����Eh����He�S���_����ϐg�#�'t;�`�~�'���S�@O�&Y }qӝMܨN��oh�7����)p[���,����,��D��7��I5��wB�C}�A"ɤF�	z�J�V�݀O"����.(&N�Qj'�a��w�$���k��g����-���aV��]ɓ/��=��VL�.��H_���2�!�#S�,@-�����%���p��|RI�J��@�r�6)�#�돈�/�Cq�e{���u�rz������OȾ�mK]�
c�+�[�f�������8��,߼�;�aZ{F�d��f�i#�%�Ԛ)>�>DH�%�$��~���ՌD�e�y�h"2Q�|ծ��M�39e�w5��M�֡�=�DՃ`�.ʏ�绱?���KF���{��ڲh����k��m<P���J	�>����'ǁd~�] G�#I�Ǳn��W�Khq_I���o��Y\*[�O��/�8��
�ϡlW����*�#9��ɽ[V�^CMe����魊�g�G6���r��E�}��6�h���Ƴ���\���T����F��{;�Rn�34˾J�i5�=MmԠ%��Ot�N��p�hv)hmI����_���z�%?t)�����CwH@���i�ً��l�W2�y�l�'�,�{xBI�<m$Uس���nI��L؞麃3:��ѣ5�M����27��IG<x&�8ٍ�a�Wti���_�IT���]y_�ŵj��;"k�بoR��4<�}�"7w�9�w[}4��M�L?3���5��@�ߎ}20ߚ��>3��0��ׅ}x�X�A6u�e�'�6��C�Jz��dW�bum�'[�J3�B�P=�#K�[�9C�B�P]k:s?�}0d;XnD?߅k�u�EՂ�@�r�6)pZw7k��s.ŧω;����r��}�ai�b)]���y\N	��7��(��AG뭨��|c�s�K� D��<�EB��HA�Frb��u�x'#�����!{O}c_~������C7��M����E�2�ӝ��.ݱ�F���]�0�Eb��7�>�Vzh���;����/�="4FM���<��PqY)���Dq��ס:�V*�����)��Kd�vKt=+�G�(�'s�3Z����|#Or�L��x+
�]���j�"J�hƒf'�$�@ܰ�gW�X��&'Cbz�m2sGj+��>�8�zu�4�O?W���������� ����#�P?ܧ�$?�Mb/��$���J9j�W���0�g��C�K�/�r�i~��}��?������s��QD��;D<W~���M_o���ʧ�+���o�~>?	a|����h�������v��!?�k��?�m�&¼Z}��/q�@�{�K�/G�eξ��������ߔ��`��V�I B�.2:M8Y&����8,�	n4�@�$)�:�=j�'��������kZ>k������
�)�}�h�������J�O��[����ߌ����o�b�۷t���I?��ڞ�s։V�$֞e�&TQ�#C p���0 �<[�(����I3�)�w��>��뜯��;�*��%%Y_���l���}�۷����_~Н��ٿ/�����N�u�y��W��iͬ�IWi����J����|��g��{J��{��Nw��8������c��W���Fҷ�z����>}�&ǿ�~�dE(='���t��i�|O��Ƈ�3kI[Ͷ�Z�K[<J;��X�}?-����|�>�~S_ׅ����� ˞�e۟<y���1�`�W��I׸A�׼�\$p��!n�LF�zL�p� @!Ⱥl+�4�(|5��{u.q9��)c�W�Ǵ�>}����_����v���9������S��[�~_o��-Y�L�_�������y|�||��H)1�C	) �G��ΜZ��2��|E�$��x_l���op��'x֜���&9�7�ZU�����4�7�iO�~x8xy}O7�8O�����q9�h(��������N8����6��Aw�P�)�dW�UD�d��,ʰ��@�g��������%��?�^7�����O�v;�W��
'�P7��~�?���}_�y�W���o�J���-��?Y �@�~}5}a~鍏�PO�XW����C�}o������0�mKe���@}6 >�@�>�O��/)��T�$�@�>����f��>�l'�%Q��RILch�D�x�R��pC��a�w
e��ۏ���x���\n^�v��0��kO;γ%I�6�����`
Uj�M;8^�$��Qi���7��!aʵp���(uݯk���n�?w�s����U;qQ��]�ӓ�wΧ�s8�&D�y&�y~K��B��qg[�l��yuJݠv�d�/O^�ӊ"���a�����s�p�_N��{ `PK�m}J�D:��=�~�#qH&�����x�����Q�A�B;D�Rj_���*O>�6d�r̶|=��v�Wg$)ۄ�Z%���y��>�ܺ��{$2	���ioqjM��s��V�`@x�wg z[C�_5�$�w�1c�F�o}�U�ٵ0,��W$��s	O+��5��H����"d3����j�w�]��}�u^L�v��海���Ѽ.�8��R�m�E����6d���L����G���iNq|�p��-�2C�p+.�*O=�u����e[����#(��]]y�W�Y�V�j��]�r���Cs�rr�b�n7<A|�-4L�5eTV[7`}%���<�mN��5-��ڤ�WO���¥�\�;%�5���>w��ff����Mw�
.X"��ZҰmk��NSl�����'G/�@Pk�^�.�Q�i��	�sRIPk��2���X;p+���F�)�
,��d[��gs��vY�b�*e쇭��W�<C:���E��iZ6�Ax�,s������3{��b���E��@������|/��(��0
��0��M�;Ņ��=_W�B��w���S2�*p�c�y�6S���H��V�!��	�g�yw���}Wf#S���Yv��Y�?�a4Ƒ�Y�e�&�a�4�%�g5���F*F��Q��2[!I��Nn���D9�%!�^)n�q�:<��6st�;�ğ�@�����󡅜	#"^�(���grX	7�c�!�� ��c[\:>-���� GF���|���^n�)��̢e���x��xC
D��g�?��/��u����t�9�����/��~>{�^5�6�%Q��4�5S��n�s�/�y�Y�҃R�v��N�̵�t�^�\s�4=�G��w�K�}�fF�=	�B�N:Rfw`�u�xbϤц�h�B0a�in�c�45�0i��+��/�P�V����fF���y��K��=�`�C/��dā�N��cz���ɣfڦk)tY6]��NG@�g��
�Ɓ	���dM6N=�b�&'F�8���ܢ*�N�v�bׂIc*��˪�/�?]�=dƝ�ҫ߭�7ELzf�z��UOv4�2O�,���Z����h�qP���ƚ=��&��V��K	~�:��A2L���yi�w�}�+bm����]�5�*-U��K�W,r,׭�19. ű���,��=3XfF���^}����2�ƛh�+�,���В�ĕ�a���E6��`�����_z4�&�Բ���c�G��|�T��ts�Bzo|����6����F��,�b��x�늭��fh6YH$�d�VFN
�<���I�T�L�Q�c�T"��om.p���M������Q�\Vm����P�6�$z[E��r�s�re�6z5|ɝ�����l����D�:(���xCzǜ+�u|�_8�c��U>�BtG��N����,�hK��T\`�Z��B�k���GL"y..M�mC��|�y1��p�z����Z�S��_�n}[c��ސ���A�;?`8*{�f��^�Ac�3�׾whE�.�wJ'~Q�f�j�2�|z���A䎩
�H�_�+��բ[�N��k7�����I�؜HE�v֫���ת{�-M���G��޷��T-� �ɘ�����������Y\�+�/1��_�ǐ�4kD1��Ɗ��-pXח�B9g�.��V��Q�[���WD�!�5�����!��Xgg�%SJa��1����+��"�.F��x"-c;6��-UL�=Y~��.��joP x���%d��1�+����Pi��dL���%��E�S�$ 5������_�u�9�:�� �R ( ��g���?8%}��_��Q?0�{����Y�&P��Md�0��X��G��adM���~�n��c���v��?�o�3�y���ϟ1�Iڟ?XmS��q�B�+�'>>�sž�0�&��|�?���_\jg[��Zq���/7Z��{k�u^������:��~	�oΞ8<���߁}��~x�f�[��T�&�.�a���_V�zF9?���񁟄c儑��6��>��wn�����b��kH����m����=�3�ZU����1���<��\��q���gƩͣi�y�O�Ǯ~|�|6ǋ��v�=���k�be�������~�㽪y���y����|��k�Sq���ƽ�^�i���&=u��3�������|�t�||q�e5
̌��$��<��sHٱ_���5ag�ֵ���v��
��^����|=�X{R��{�����M�y�W�^�#F�E~m�����2�/W�oo)��w�6����Z_>���v����3�""�e����z��d�R��a�"�ύ�;��u�#=b�G��y���q���^��e^��Ͽ��7l�^�{ˏ�W���ޯf����m�D��g�>G�TV�i�mD�����c���� G�GP���'�ᡢ���Y�	J�	�y|�;�x�����<���+ ?[���B~�{n��>�	%H��gr�g�4�Y^u��o����(��ξ�S1�s����t��n�b~ʜ���9,ʝW7k�j�k�����i�T�k/�hN �ۙ�O�F�v���ʐ���*�K����쮚���x(ࣧ痉�p�X�ퟜ�6r�tS�*/36z*�*��X�OA�B7q
�5ms�:;:��M��Ԓ�5���R��x�%�$-�UۨNC;V�nV��x�B�9���Z2aT������	�	�Dm�N����:�SB�B]�o_p�c�M,k.�\�r�+��K�V��$��ͩX�U�j�;<v��@Я��Kk��.w��fm�c}�l�:��n�7��Mq�/v�[`s"ca�����+l��r3�;-+����ئn���x^>*�r��.;@B��ӵs��!N7mN�um���;6�Zs�'nČ��-�ۙ̂Ni�Op�f���ۙ���T��r!�q<�ͳ[�劣vF����2������KS艾<�S �n�F<�=.LM�g8��̬ͭ���q]m+&��sy������Y�%U!e�髥�����%'�,TPR77#z�;�q�җ�	�ț�Og��0��ki<����w�vd�7u�zJ��u%]4��>�Z�$j>��z�u��:mO�Ӵ� �� -�؊����=w3��9Mҹ��^�Jv����a���gI��}��WS��pN�r��
n�"��EXQ�.s���sRJܝ�8�<I0B���*��2��j��w.p�oh/o	���Mfګ�ja-VN�vt�ٞ�ۀv�]7�z�����̹� 1p:����M��Q
��ܼ�۫ч�����Y�����҃�����f�/��������R(;s�s��7H�}ہ�ԧK��D��$,i���FN&�\SSR�&�pi���2��,A�=gZ��ܩ�b��Y���	A���Z#wTelė1����z��Ǐb\R쪌�흠���J*3!\]V&5�򢮱wd�Je.9�q�$�{��\��:6+8�kW��l]��ۚ.(�kd�\���#�&�b�����%�3˅�Y����&⊜0��0���R0���Oic�� Q���+��A��nq��c,�*;N� 9����k0+�nY�49o^��+��>���A�x3m���9G��#x�
����ۛ��o��- ٱ���TF�{����cvpt��h��u���43��C�\Z��P�ye��c9�X��T�nB�c��jy3�դcf�S�������l`5Vy[�y׺�Z�rzf1Y1�#0|8MEVpVG`��U�����(����k�~jDwG8S8$h����܆�\�Q��p���R�"���e�)��bD'���yBX=�\�xkr���m�4�sx��əU�u^g]��&7 ���(�
���x���*.pyߣ���5F����5���cO��b��5�i����&#�D�a��y��
�}pg�B�T���4�����^8��w8x^�M=l���gQ�����.rb�8���Y�T+Q=ϯ3�nI�/w\��-ӝ�[�  UF�=wutw��Y��!� �Egj9����;#Pw��B����8��)j�(UT�w?Q�ݝә������1�j%�ZP��=��^E����G'�e	�f�c���3�V�%���U��hf��+7ݞ��fMK.���T��P���sw��\+٣�n+�kovj���錘9��s�#�n��7�
��,� �;�Fd���2��]���e���s���j�ڹ�D�y�'��N���z�\)�3��.R������.jEu,osJ&�:�����������,��/���ʻ�����d!�� q��r�^&�)��\�u*p:R��PE��d�U�3�q�j-����SBZʚ�rX�n���S��B{]jgT8�&
�1!����9�`�w��猊�Y���ù�f�fo(.u��pY�ŵ�^ኳ� �r��1uc^F�6FLA��\�dm��]�O9�h;elެK�PJ2�^K��ߑ��^�I�p�}�Wy`�b��I�'�f2�y;bA�q�t
�[R�]���P�n4'����zxe풪��Y�Y�F�+,f���q���#de[b7Z`�ڝa̵@��mN��;׽]g/c/o׺�)$�0�M���}ef)R%Ul�d�H�cFհhӊ���jIp��^�*�i��][�/G	���b�
j7�댫1��[�J��J0�p��wT�;���ܼ�r.���b��z�~^٘��T�a
�Lg���4�n�}B'p�G]������^��|o]tT,9����^��ZB�7�uޒHs�[؁=6�1�zw���n�ܺ���Fa�`��E���=��:�z�����j��m�8���@��!N���y�-��Fs2%���u�J���9���Fs�U��D�H�������b���gW\V�I'�'�V�n�9P)�v�ik>7۽5�"�u�cf����k�e̻&�ZY��Ou�F'y�٭g��P��+��\O-���m�sPH���#��o6f�±#����As6���]�GGl�O����1��Wb��X�>���Qη�ܟ��ݨ\��	��vj��,J���cu����ʒ/��F1���C�a�p;�Y��7{V�b�����W���&�j)�ڱp<*0����U�TR��p+��7qW�	�ŏ&���w&��q�9�9׊�r/�`]F1'*�����Vj3N�yW��R��N[=*��׶r�Mf���-Ft��e��Y1�K�����A�|-vc����Mƫ�����W=�{E�[R-�Jv�D��P�Ln9��W�i����:?WLl�&���g]�Y0�)9N�T���)4��wU���"�=q�f/i�'���ءwj��<���Tn�/2�4ˍ&�ټ����ޜ����*�gw�[FyAT8�a�ϴVl! �V�փ�V�m�TQ�|�el��v��/-(�$��b�D�sQ�p;!���B�ԩ9�'���9�8`��|6���3��P�����`_u�m�a�&1�5��6�j�[H���b��v0`(�Z�G\�d]_�"�=j*�L�xgnt]�nͲ#L��W(�R�G�/Y����\�;r�y�EK�b��U�=t�wn�o���Y;�1=�����V�vfS��X�f`��ȷ�t'�_�2�r����sưF�YS��O���z�zbX�h���*�.boX˪��8�ܢ�lD���g���P궮2o�=SdE��Sa��}�	�FЍ��Nd�t�sQTP��'v)� �f%z�Q��fk���V�ܸ�����kSU�<�{d���Ѷ��Cp���&D� �ͺ�u�&����V_.���w3rj2�F��W[Kj��uNc;�1u&��iND�Jܼ�3�5��.�"y� "i�J���m�������k7=
Qޭt���%�'�:H˦ ��T=Y �p��7�<��<�,��SA��/�7+UWV�xؽ�x#"�\]����z��DF�J��ڃ�9�\�F�E��{��ji|niw���z�YɱA4�<�t�s�l��4��Q��ܘ���cb,�d���MK췙J�p�u��L���3�2%���g&M��ϑ��ng�T�Nr�����8��܅k왾�xv�/o��\�9̎���u����oNQ���T�����:MTjF�i���{�^��n��F8�)t��ʹ��|9 �v�gqȧ	�"�f;���-Z5L����\��G��=<�c[���
�c�cٵUX��S(S^ڰɿ��hW>������6fPȰ{��ˬ̸�Yл�w+��&��Bb���F*ڎ�֭��X�;5هg�
���Lb���*�U�Gd]�N׆z��׼��JY�~�5�Z�:�5w�Y�qFc�2������n�An�Á�չm��Opk/$ہ��؈o�O�S�v�W���VƁ���\'�)+ �N�>u�\ogs��ٝ��w��9(��1=�뗛�e�ݭ�w�\��,r�<[��������cpF��,H�#+�F}5�L�4�F.���]]�F@����æ�s["3s;jS�Υa�m@�yO���]Ob�U��]c�_��~&k���Գ�Z��*�<�|7Ը�[UE�,��/��N�5x�d1#]Ҝ��p�F�4����u���F������s�+�wݫ\�otI��7�����!&�J[.jVK:i�N�\u�
��9��/)��ں���A��g�j����W{�"�u=�3���Պmu�����m�\�=��s��2B��jl�Yi�޳�9t]�׏��ݎ*w(�y$��K{��gV��QG�sQ�<�_c���}�11R�ފ��_T"bLk�2��A],�h=ܳnՋ�.il��v�n�9�wd+�燎b�b�3�����O=!�5 �۶�f皪}��]Z�}�*��#iK�u����^W[��Q�SW��s�������n���ʫ��:��[���Nu���|�� %3���!l:�ܮ앀�f^�_lζ�u\�t2��Y�9���N���HA��7�� zҁ��+�n�q�-Аx@��&m�j��9�[/6E]d�i�9����	���B����iV�d��݌ޭ��3k$=E�����C�@	��^�#k��V9�����Q����*C
Z�sU�� U���bo�2�PP'��iq����V5��#��4#��!ɆX!�{Qu�a�A��a�;�a�Ma0��ݒv�-P3**�W���+k�����7Q�ĺbP��J;,.죷��9�Y�����tC��4����p(��U���3%f�|�B�ܴ����g�77I��͌Q�/�賙��66�W��rO�8ۻ{³��Q(�2�E�����*r���銹���� ȯ�GN!���qC��W_Lƚ��j3x�����=���;%�^d�	�F�]�:1�W��vB��R�o=-�Mn�&�1�^h�n�\��<%���v�-&�ʺ��r��h�=ax�4��n���'�9��ں�&��.#�DN�{%I�`]�Á���9��ٻY���W[w�2���@���.:c.��jpU�ǝW�EV�4`��0WX$�=��}1����������;9�����BIQ��'b�k#T�60*�L�3����E�:e���P��btV���lL�P�u���ĽѪ� {�\=�۲����s;4ʁ�c�wkhm����U�8���F�cIʥ7 ����|����0H
׷�9m���sKg Of�٨�AS	�U8�`	���w�����{��մ��wP����c�ݳy���!�5�q�ڛ7fPa����/�J��fΉ�'�,��V�����~�y�c�)�'pk����5D�(�Or^l�f���':W*��O��n�����Pz�Q,����b���:�cy�����B�EIQ�BJۖ���P�!ᒋR��������.�9z�6#.n26��&����t���{��2��5�1vVntp�y4�u�BC|���uP�=��36�uXe�&��&��f5�9\�y��OW�ն�f�\�-��L&�m�8�Mɥ�+,��PDe*v�Z�:��օn�v�o�2��Q�p�U|#\���~�wzoO��D���wAd�7�'�_����z��iM���ʺ�f YV)M��sC�fsz�,�պ_:�E�s�%�ɺ�v�j�QY��ƒ�{�,B̀!�v�̰�c�QاI���I�S���M��4u�2l��Ǻ�Ud�uYC������P��ٶ*�Z�s{�A�L"u(ͩ�
(�ȫf2���ӱ}a�z#4}]P$����Yک�=t�m-�;�ۗ��ļ���L^���N0(��Ӂʎ��٧���>X�W*t�v�szڤ3n����GnA��]!ul*�nTow��%nK�q[��j�:�#!�:\��޵}}S-�ƹ�:�vm��;0�[��͹u6��Ov��M�
��Yݗwy���uq�L!sYƔt]v���lV�ۋ��F��N���6�g���v��3Unb�΃��5��s��I�fS�\iNO%$�Y�ԡ\�*��Q�'0:���K��2{0����E�	������O��;�yV�S3��+�.���8\jH�V=����:IJOl^v���&�mf����ڡ�Q}RI�kc��ЙV��n��4f엝��}�I����}���z�7WG[{����8�9�l1b�OYU�R.o#�O\��e:݃�	�[[11�LU�1�n6��8�ײ��D�^eݪ�����)ޡ����GwK$Y��WR�la�=�y��pc�'��a��5-���-ˈ�講��H�t��[��.'W:Uي2�R:�T����Dj��Yu��9[.;cV�>��;'p@�����=�d�>j�M��8븵22Ůw,��4j`Z��_M,R���J��\��;j��\��P8Mb�̨���	پ�Ó=jz�e�ϭ*��R�@p~y�c�Lm��@�����-�t�БOI�r��K�R�z����X��hm����ջ�\��P�LWVe
�!��pq)5��H�U�,��&������� ��j��ΨhH�w���s�]WZ}��[V�隝ꬫ���w��Jq����)d%���n��������D��5q`H
0�zq��������3{��E�Q�O([Wpa���N旤;�D*u���j�^ܷ�'��*�%��$v�����������c����nkH�-�VF`Ef�N9�yǲA����뤠X,�ՠ��sTc�WwNot���GmF	�bR�l/���J3\*�L�nΞJ�
o6&�_;��F�M췈�Vz�`�j,��i"��C�m��UR^���/N`����E���i_=��86��c���=��V�v�sI��O�ިnF[��C����|�#�Y4|�n���-Q�v��-����{��{�s����u;T/R��YrN��R�ᦳ'UIy[+X4G(}����6+:�*؅�����lj�xIٷ����Cr��;E����[��.u^��p	���FwS�o��ŗ}z�#`���uH@�3�QG�oI�VVt�����7o�S.[.�[�����s\��h�*:,C��CW\�d�r^��
7Des�p�����@���WZ<����<���36+�������!��@F϶_xQ��l�Ú+{���.%Ui�L��n�vd�x!]F����,Dnf^̍�;0,q��e���˰��N���R�CX����#������d�X��5!��vH$��nXc[�����q"mk��(=��gX��^8�Tr�M-���<VCԵŠ�9Ȝ�-�k�+�'ˉ��=�b�j����/C�2+�69e�/\�W�y��3�C;�+V���Y�ا��&%�);;�l��}��a��sT������QWvn3*v�WJ|��]^�MuL"�Ev���Γ�BB7^�	��KS2�qUV;���!\��;�CZ�(V��q�8H&�����xf���;�e���t&�[�7Fc
:�7��,��#�L�"i,�-�{���5�l��/ Wa0�J����@�T�]GL�yF���<����st[��o"�]�Q=Wӂ�<�V2���6*PM��o��禣*���dX܎t��#G,	��n�rD��24��3��s,�i�{Uz�]�fެz.��ݑ;N�G;X&T�B����rd&��'!�.GUt�=�/��쇤�[�W<����2�QG��#�7���R��U�c7'h�2D�{��}st��e�G����b�z	k��3�6�N�Э�Sdd�����6��#e���\�\�<�7%�d��uh(�W}�]��UҬ�_�`cs�)mӉY��qӫ�/��I>�2��:���k#kpm��]�Fm�ƻ��փ(Taz׶�hK���uR�㳗Ps���\G���yǫ��[TT��.�DfbΑP�JsTH�mQ�s@�'X�&��&�Zɜ�-�����7��6n�8n����tJ��֓;�D9�D\�sx�<�a�M�(/i܅�/9�ٜwm�1	��J��f5EȒ�U�����;���[�zʪZ��"H�Vi�%��Ȼ䦌k���*F]�o�T�����jN��ɅJ��)�ѲL�0�;�j�-J�7�KQ��o/,����
�w��Xь��	�2dvW2�$_6��	%		0����3&�kǷ3��2�f"�&��'�p��[{ܢ�ɹ��ᯟE䖊�g]�����^�r�.�kNᎬ���}�fn0��ڥ��������S���xuF>u[�.��2�t!cfj��$��f&�5.MeZw{6�&&�D�Q�h�̋��]^���	��P�8���+o{̨@��4>yS7Z*�W3��-V�D��s74��E)�S�U ��8�{;���63�\n����(��d��}+������c;����8rν껬T�8F�q��O�a'b�=�m�N�ІUWiZ6�Ύ%^���ƦD����<'��.��f�op��$,����]�2�*�w��K��Vm
�(�j���8Gj/��7{J�7"^�;j�T��`����udPU1qO��{�˸݅Ո�mέۊ3N�brw��MZ0��,0~jo^����T*/�s��Q[x�Q�L}�׊-��A53F��I�TJL՗�/*��B�o���RviE��.��Ef�c7�]-��.F�������3�uEe��NZ���VV=��K�;�l�Ǟ,�ӱ�5L�����Θʪ1&�gLw
W3R�L �ͼ����f��X�b�gDU���nzo��ڲc���NN�jfM`CY�v��9�;gT��;
hBv��oLb�́�a�][8.��7��q��q&��=��87ɩ���������^Wu���y{Nv�{KM�����n�:J1k����Tg��TYhL��[��e�aڪ8{��'e��W9��9CfNMQ���qͮ��ҭP�KU���m�ޱT�gO���3��F-�s�*��lاV5t�ƞ��OE�����:t5}i�0N��Es�۵��*TKbs��}uS*��+c/:�����̽ڪ0,�S�$��Xv�t�LV�koH�����F���V�g8�=�jb���bjTGBsJ+�lD�/��T��j��$勬��Q7��V����f��;%���Sӊ�So���N�Q�1�Zڌ�ѸH���&t�,|�7��H�;��#9�3.�p]oe�e��C��W,��sA�[׵91cQ��2��[�������/�n�q��F��-�ڳwe�9�@-�v]h�ZF�u4@[o�䝮��;�yY�\w*��X�W17���2��@�h�f�3t�躛B�*h��])��P�8�꩸̑j�x���{���Sd�f��@]��4�i�3�N1���wTE��sqQ���O��v7vn���@��k)h=����"��]=P4o\�u��7)����T,.� |e��}��e�W᪠vp�V;�L�'VgF���>��)��,� ���˝N�M��;Ҋ٩��T[7hȮ�W�JYWd�}�*r͢�xv׉��1h=�.�j�dl�`A��	8-�b����;F&��̢�.��p�.�@W-�R�%K,cc�BÉa6��u[���H�F��AU��r��:U]�N�e�����:2�&:ҫ�c�L5IKrS��_AX�(��_<�uM�페91w�f��L��nr�Z�9�YA58�̈�SSt6�L�s0#bp[5g׆�:%]Hn�I<s2\��pb�Ps �5}A�E@�7r�+���5��-e�7�f���w}�������L�G�멠K��E�&e���C2��+J6��-_W�
ݚ��W�;$']��3�Bf��$�т7&(M��n�)�3�@�5�%J�s.��6$�ٟ��73�q�ȩ���U��ս�r��l�]IЕ�G,��j�MTa�z:�Pܒ:�L��vAq7x7]�c����U��TY&4b�)�mЎ�ܒ3-s��1t���_o
Y}�99�7��=;(��M�%<3�¹D���I]!��F���J� �6&*9�����h��Ⱥz�R�V��UX�K�N,�������.���/��g�U�@{�·�6�(���j�Q�vu�NEm3Y}	(�&0gN�)���v���Qu�	Tr�u
�Ǣ���Ҍ;���Z͝tdF�6���2.̔2&�j���9c&{Ӝ�lI�B*mKꞧ]�YȦ��
��Q�ά�t����m�c���Q��3�5O�6_pԇR327�M�wN��Nl�)�n���^h�5'r��;����*��������Ƕޖ���wM֙���ڙ7�ZU��g=��p����L�5�+ ���{#N��4]j�`V�դ�VK�E��Ul&K�MX��n6*�-Ժy��5��:0:2;�3�R��bud*Ω�N�F���Lٓ3/�Z�P��
��*�M^�q�ҧ%�s���v]��$�i"ܩRV�O/s��b��f%F�]�\9�����I�����C'����fLQ��]3�We�JيY7F��k��e�k�k�P�;dG\�{7s��ɬ�z�ue94Vw�P��ycN��+���r�'=Հ��]�n
l���0J��{{��9����c"� �Һ�Y�k�Q��[���}��vМ��@��j�S A2�i�6�wv.kn���Yd�L�=o���s�j���h��T/!���	���itRe�i�o\ع�fj��9�+�xA� �"Z��&$�f��1.�n��3/���T�CIJ��lSʫzz��=�����q�bb��N[��I8!8�I3�"�T�1ڳ����j���5A&�Z^��u����sې��FY�iv����vHۡ����ٕFks:�84N�c�6+��B-���
bz��B{3Gp��B6�ùU��Z���n�sr����UL`a��tx�NVOE�AE�&��h�T��˱?׀���k��˝:�n�1ӊ���M�]�m,��(��{ݗJj^p�p�����u��t�m��B�����CRc�]�]U��_u�a������L4X��B��L�;K�XR]�C;7��`�s�6{(h����@(�оW�/yp���!�
���ԝFw3+��T[E�)�U�ngUL��g"�ܴ�����hy�r���aBʎ����]uoS�q���r�f�HU��x�q����P�Y/����wa��Nq�,R�1'����NJ��{+�<"�n����,�n��e� �Q`�\�I;�w�dw6�S�����$��Olm�A��Q����.�$��q�v;��ȭ��P���Bu�4��H�޼ѐڻ��8��LQ��UZ��찅w'w�+��މ� \v9ɫ�H���x�
�]�]�B
�Ƚ��#7b�e��G����A��_oN�s�oM��fy0��#�s�����噝���ub�_v��g;�FJ�6�7��i��֗sS �|��9{��T�Ժ}���W���X;�b�Yّي�B��S1Z�Y�#��������4h� {��+X�x��u(ѫ3K��0m�7b��V�R.$9�q��A���L���n�cx���a�������6`b�=��%�ͧ����YUP�*�'��T�a�*��8>�`���U��i>�kqjɩ�ړ�Q�7�����*C�VlNh��U��G#@^�*/$w.��~����nB=wq�OZ�=����`�T���:��^��a\m�+b�y��ᛛ�� ��;<1h-�꒶��u�w!h��{:�\�G&`Z�^�%-݌FuIQ�O�%�Mq�8�S�s�\)��܌ tt�zIu�I�ÀU�9Գ�-�ޡ��D���R=m�e���|6�s!ft�u��1wa���7�:"F�C��<�&)�v����U)�}�t��rb�mb����������'��Uu������;�c"�D���v��z�w\n�m�̸ʺ���J��yU��o����1���gV+���&���v���˫��\�9:Gd����YΣ-�N:�g�B���3���˄� �����ڌ�n��·ja/8X�t�rh̎���1�1U��O�6�+�!�3�m�������.�1Fɧ��3Um��vp9���:�a��߰����u5��,���{ʯ^.��l[��:�-�ﶜ�����v6�v����uRyuU/��w��w.�"q�Ϭ���gC�jr����w(#�)|���૕���.*j[��^^�̈́�"��PjV
�w��fێ�����d,�p�-����W1,T�����3�T)�sS�j�-U �tf���̋]'}��e��8�ߍ���&����qV.�5^�y^E:�S��d�]����wAk�)V�7d)SAIa�o���!ghlM�T�v��yئ�.�v0*:fS�/��Ż�a)�o��u��^��n���9]�[�zDl-fULpYԯ+9�5�l��,t�G(>�,�Or���ua��H�A9��w�h�I���@X��=f�8i쬋ᓎ���s9�Y�����!��W��2�Uw��ל�����۪F�s����/"l��ݛ��u۸r�v#��и� ��ؗG�%S��ҫ)�BU�
;hB` @  ����j�\ō�"6�؋4Z9��v�rL6������ܷ"��W-��\�5r�d�F�#m�&�[��1���ZG���\M ��oF��~��� }��>�����O���9���?p��\��<Y*�_\��c�T�W��g��#��,ϼ3�w|A���Β�>�2ʧ�~��aL�BIf>���U��+���߱4R�Jߩ���Gk�}���~�B���e�}��`U�dkR�U���˩J�4?���Q�)��?��:�5����F�d���^��
�߂AQ.Ty����O�Չ�q�J*H�Q��s!v�W���9����B+J�)Ԭ�˜�%^ěE|��*�jW+ws��N�y���o�{pw�@1�EO����lq1�|p��7k'a4_5G~���n�����	�(��7.����|N��tjpC�=����Җ�P��or�̑�λx,E�j�VϕK�+a��,d�U�:7��X�}W�>v�)i�7=K\���wb	�;I�VtU�UR�+��z���\��˹wڼ�~])��j��]��"��n����Hk��?P0O s�=8��a�eK̺��`dc���8s�|��z>��u<I
I�b��#ז�1�%7f�V�Ԏ�t�᛹����e�0�3£O:�^�De:5��� �Tj�X�{OM�f� ·��`���*�w����������dѥ��/�Rm�z'`�$�� ���{j<y%i�,#�̀v���ԫ�Ǩ�Ȓ*e�{*l��E�inaJ����'��숻odӭ�v#L�Wf����y�b��*�z���
������[~� �<<����\£C<­�뇟S���?Xg��'�y��}Z0R����>ߟ�Ԕ!�={;e'
<�K61��{�8Z-�a���'���{p�T�ĉ�����B+�> ?v�J�N�*��ʈ���b�.����-� �m描�Y�U�����ԇ��{'J��ϢG�L2�g�\={�S���9zfz����3X�7mug�gֽǹ
n3�]�b��vv���0D�U�k��.]�Q7q�'T+,�Hi���w����������Ӧ�����	����oV5�'���Zo}C����u�1�������#1[�Qn�-��o8>���>U�3���$i��Qs}h��i�{Վ]p�|����L���^E��B=8TB/Z�
B������:ڻ�nn�|p�xuc�nί�׬(e�ۄ_���^I�*���"rRF�R�|?+cD͚������~Jy昸0Z$G��_�3��{��P��{n�ǴM��̼
�� OI1��f1�__�-(� 2ޢ�(y$4!�:������pG c����3-7U�́��#�a�O,�����SF�^�U�$t�Dq�� 4u�/�A'�l�%"��-�r�p�ޗe:r��z�u͜���U�����Ae<\ϱ1$�����C��߲)��T�/�+�M^3R�2�Vn�u+��ZDb	f(&�%B�J�z�؋��հ���pO���U�7�!q���F��g&E5��p��JsB�ί G����z�L��(��ùb�>F{p�9��?.�=�+��Wϯ�Z����E~�������6� =�����ގ$ޱb�3��/��E�
�i�`�6.%��)ݳ��!��ண��^��H�bI�H0�].�O1�w���a�~��z�r��]���1�k�%p˃����G'��#���do�օ.w���|X(��5�X��%�`��!4����q�H��D���Oe����(�H��T�c����	Pv�� &k�z�aVfU��rqr��zd�<b��mR(*�������z)��|Q�:�я}{����p��RF5�~&6��FL�J!���JM�g���FQj�W���RW�:Z��c��v)�^�>-���k�BMq��B��6��<�fw�u^���m`�:e��O��S_���ܢ�ޱ��_��%]F`]�[������ ���J,�wn�
+�m�S�ǯe�!�!/{�zi[�SZEޣ��;R�xw_���({��~�yV{�h��R=��Dܞ����$BsKZ��'^]nT�����a��.�INzP��Ed/vIQ���5���U�n�0��vJ^L��-�X�; ��C$��ܿa�X��17X��?<qs#�$�WRڊ��R�29/GtPk�0���;I<�7��&�	�kP�\E��Ř=+p����szB��q����L�Ƌc�|߇X��X)GW���'x���2>P��Џ�}�ݯJ���jA��:�����L�Wd�Ջ�}_O�>�I$���z�?�8Q@Oo�A��#����@xƟ�?o�}��07���cl���I&z_ٿ�_��H�PQ��]��Ï8�8Y{R3�=���$�R�6g:=t��z�i6��ˋ��)�n_�k?����>ԝ0���������uꖰ�+,�}��E!��Q�1��ds9߷f�oTǟ��{�<Vӓ�c�N�c� �7�|��=�����od��E���ھώ��i9�9��x��^�5��JTޒ�ѫ���Gi��ǅ��W��v��Mz-7ǭ`�T/x�{u�_[�]|zy�<�#�#kGd�I���_k޾�	���e��׉��o��p�o${O�iO��v������խE-[�T ���6����'�
�����j�U�L5+^-�Z�bm�꺟~x���6{��ϧ�%=/�h�:�u������2h��27�.5�TY��ݔ���3�L[Y���������T�ǥF����WO�l���'����f��ۦ�Oy{{_�n��|X-���jǊ~�!G� C��P�1� `����7�~�����_g�z�.5���P�
�x��xO�{�����C�r1���F^������������D�k��������?)��G�R�E�����'��U�?FL�)\'q�2p?^�ѯ�^�����,���~���D'�Ui��}>�a�ڞ�U���q?q)�����[$ ��~Ӊ�~Ƌ�r�����<���B�$=�O쬌J�Y����ӏo;]g�КtH��V�wP��l�!��][�m��}�a������D�Mb�sF�,�DK��"�p���u�s4VO��no"�I���z����`� i��[ޱ���i�?��S[�x�mnU�ֲ��=t�|�.�S�-��>������e��\�����mZ��2�l���.p�K������)!��G#j����`-��d8�VFG�@OZ�;�G�^
y3������|2�-�ڄ���+�s�����Q}3�s>XT���%�(����,yw�T��2	���h��&>���tr�R�?T���]q��o
����H�Ʋ0"�kyE�I%���@׳���Y��я��J�h����Q�~��~pKHq�:��
֣��O� \��pI�m�%�Ԛ8�CA����xg3��U��^Px�ܧ<�h~ǣ�A%�������NW[(S-�	�m�P֒��TL��]�PSgM���GL�.N���~JQ�X]m~#�hF������M��fi����쐦�<syY?L���4E�{�cb����M�4H�y���&;]|���q�j^��_^�#7viǧ�Lda��Hv%�,�╩
/���]�g,��o�X�*�|=?:��w�*hV/Z�����*|�]�-1��zF�z��b��y��;w�o�Ӿ�߬ʈ��-����a@R�L��>�B1o�\Q�z����Z�T��n�����0=����h��X��o�m�*��${z'�]h���y����&ņc����w��ݨZ�8*��P�b�p���T�`����_�n��.1�?�I,�L�.�:!��Q=3`��w��c�U�W~�
�zꔘ���^5M�2`4�6zm�5{�^#f�YU����#A����{鍸��.���g�� �i<�9�]!�S���ᥚ6Z�¨���Ksq�?!y�n7�ėO!K���h�V� �����=*�}�m��@�t��z�EO��Z�M֒�Gp�E��щ=ό�sf3+"Xq=Er�3{�����_��	TLݶ����7E(�E�w����d��ד��3tS ؽ5r����ߜ�v�|�q�#O^�k+=�O e?��,���ݦ���܎"���<#P ~Ga|g�k;PcĚZ�[^�ܚ�=ٶ�
¹KJ��h�l[N�F=n�hzP�j_�����酴��17Ћ��A�4�-�rG|��b"oZP��(m���ER�2��~M��Ϟ�*o�v"M��ˑP mWԂr$�d�3��r�-�4�U�svׅpنw������.�Zem@qFk�bTIy����M���5�6�;����`��ʂ�]8ʀ���^�wݮ��Ii	���b��LSq�Z�1[R���.j�X%��_p.v@��|\���PD��_=,A�]ѕ+̗��)��@#Dx�,���/w�fA�V�%���¬G���.4i�N~�!'O�M�I�]�%ã��E:��f%�e�h�J>�Ǟִ�E�f�8��|b����O�u�.U=�q΢s�����l�	��ȓ�yn��
�d�)��5�6ٴ0���ɳ=�<��"��[�x��u�\�wꦍ�]:1�����ħ�J���M���ԥ��NZ%odٵ�`�B��������o��I��%�bh9q������Z����Qr�ي�,�f�j!�l�P���b���7�C�Ҭ����&�y��}d�4Ƒ���!�KG�V!ӆi}ԫw�'8 �S
φE��l%��>���a4r�d�ԇM��[�s�mM�㏑��Ȇ��s̫��?wN��IfF�y:~��S�#��avncY��o�M������@�ڒ��60{`�| ��
�oG�I����~?��8�̟5(��ڶ�e����u̬ �0���w_�揄�p�(�ߍ*����� tP-Wuw`>�.f
��N�TU<��hl�V|������+��u4u�Q�4wl{�<>y��*:Ed�׎���_�׽��U͹�:S���=77B��n�]W�|�p�R�}m �ADǕ�/�|X}�i��S����H=�}>��}>��H�,=�Do�'��>���H}��XA�LT�
C�H戟�L߸g�8��4�k��ay���n�35�֠ӭV7�J�]�;�(�C������y^�٦(���T���z������U�;�7�}V���;��߹H��O�Ίd��D�i��x�ﶢ/Ů;RW�D���΄��Jh����,���O�3IR��x\�ݶ�+�����0��[KK}Q����3�*��.���s<����&9�j�L���{q��C�����F���zp4*/ߎG9�D�Q7h��F\L˹�H�����Z�wTJ�<�;6$���XJ�i�f�d��{���w9A���zK�J��l�*���'�y��=���h��|���]׻��X�;wJgiH���ۥ�q߃�:���m�z��CU=�aJ޴��[�nki��w8�7��@�"�3���@�D�`?S�~W��'s����p;T�}�����ؓ0�&�f"$��(���=3�׋s>�9��?L���":�.�>=>P��*͝kܮH��Mk%(�Eڋ�u�UJ"�YU_�Sx��^,�9�o%�n�-��pV�;�4�+�')I�J�R�cEB�x慁��f�N�=v�;Cg���!36�FZ�x�U���1y�ՅW|Lo�F��s[�ʱ�V����q�����㳬@Z^O��6D��Y̷gZF�Jʡ���{9��2T������Eb���"�7C�Q�OT�앣%�R��xUvh��-N��d%�;�2�;�x�y��y)�S*�9��j^I�����1��!���;b��@����B����D�J��<����'�������W��ƈrL"*H�%�IReU%�	�IA�ID @  !�=�'�}�����$�~m3Uk�����ك�06��e�Z,�D���C,	fhUJH�E"se�Zy�h��ւ�Ol�sUy��{�XH��M�u�s�ģ\��:咸�����j�vȌ�g��_	т���5��Y��*�R[l�ɛ��I��FIk8����Y�Ix�[ �A���K�*�sH���IE��[+K	�5�yJ(1&�p�*"���a�"h���,�f�h)�r�˴P�0�$���c�L�U�c1WIQ%ɚ��L2�`�uQ  `�,��O�����O����_E���yJq���d� }�_�~ϼ��>�D����J�*�MR��2b5*5hBEq�j/':��Y�3
�V�b`H\$���45�WNron��U����޸�<;�f���S9�e�l�$f�+6�!+8o��uun&UJ��
u �}Z8	ͨ�D� � ���"c@���S��7�G�}4�+�Bp5L>#�t��v{�;ȁ �dM);`���,ᕢ��1f`��Cp*i}^��c|X�5�;�w�'!>>W�}`��!�O�{�>b =���M5�o��u6��]	��}wݷڱU��=!g���OI?	9���@��ȩ�&��L?<�:�����ːa�D��'K/��
�Y�\�ё�!I�p��r�3���~��b����D�����1�ې�tE��wӤ�������ĭk
�$�K*��.�i�꛻>mX��P��a�.�"��-��M�q�ѭ�B��{�,KDd���A �tA���H�����G*�؏��0-����2~�(�i�4��@=�IJ���ԛU���ӂ`�r�k�����b�v7b��e.	��9�,A l@�_��;:oDSr�A�f*�GMȳv��h�K]��ED��a�e��Fz�`(DEH��֍�����W�\�ʏ�=�a|�$I��٘)�W�k$��5�]dбZ�%eYSU[7I0��4R>R˄���d���p��EQUSH��Q:>e\���:�f��B�(,�*C3+�D�CQ�J"+$
O4f:d �*DY!2GTD��ϑ]���c��5S
��b����T�7�H��v@��I�TB�u8k���	4�j#�B�5ak!���(Un����!�z	�'Jʌ�`���]
�� 5ݩy�UY	(bBeZJ)<R5�H�w�%�4u�FHP�U�hLU'��ngZ�)�� ��J
�nU'4��̬��so�^Af76v�Ey1B�$N�p8�5�|�r���E�!A�ÅS0�(Q[��Iu��Fr���P��6��bmu�����3��i��H�E��	�ԡ�`�.�;P`q�K%L^W1P�=y��D�I$`��������q��l.S�Ad�İ#diە�ȚY!�����3 EH]T"�섪�V�h �$f�A&���fY""�j������RJ�n/��Q�]Jɔ�@j�uz���*������\'��kv���s�W�-AU"E
��YY�!����!UbU�3%QQU�d	S��"lFH��\���R{*�]��S����l?��k{�qTt�&�Vw�����x��x!=�B��W�/�;!�¹��
?������>�;1)
�k�*�A��Y��QaQU���7���H��LUh�q��"�#�zZ^i�8Vk�HV3�9�I;�gw�����\_�ck\���FEp�D4"i��Q�W�R���S���!M"2M�D�TL�4��t��
9�d�4+�"X����%��(d�c�QP�ZVP"�� ��a�z�qp rRvEA����N����kEՑ읉���/��3[�0��U�z��%B; &-����{�.
d`!t@ql��2(L"?�3���8J.�	i�X`����DO�L�K�K0YU�!�-"df,��d�О�ӧe�:�޺��S*H��T����7Jx8aE�d¯���
_���x��#����Es+��I91.�	$���
��r��~��0X���� ���K��6���H'pa�TGs�e���r��6\Wf�>d�4�����(�K���#e�!��o+�a/Z�Y�<+Q�Q'X-ȼ�L���r�7��*Ȑ�uS�[Ƒx�3��g ��BA��1�B���n%�Cf�aP�C�%F�� m��p6�n��J����9�0Fep����UA#'
NN��I�EfP˿ѹ�b�f��ة�!)9�r�D��3d���\b�ڈ׹����%s6��IiS�l��bp9�)��T１!fY�Bc=���o]Rx''ɍzg��5i�Jt��6�j�v��<�Y$�O��$�*��ķ���u��)��0�b��Bd.ګ��b<��/'����V�6S��|r:i˪$Wo��l�)���â=d�fSJUV>;�g�m�LN*F��{�8�S<P,�&���bP��R#Q
*P�D(�����1�k@�u^H�rf
 <�m��|��K�������G:����d�7��v�w&�b�:+�ڊ���m[f*A����;�
�M���+�N���ʹB���#;/"�۔�R)����5�j�����|8A��1Y��e!�!��[TF�^�؜�2��|�r��8,GM��]^ݍ��AWT���  ?��O�q^��am�p/5�
1��(D��(�AD��(�R3�z�"bn���v�bZ��tJ�`)25VӠ@N]F�ȝM��"�a�EQ��I�69�f]�u��)��p��� ��"\p���-vY��Y+�LF���QF�-k�h�R��`���p�u@�����EL)}��i�>��]�=�I�%�[0ykWziY�x��1G��"��rV�����ّc�4�򩬼.Mپ�֧c2�r���<N0�S`�e�6���nB"$���%���$Ż�嗱��% BH'.�&�G�Y_�Z7I�c�BW9R�X��
B
K��xWWxV�z�j�K� b�%1��e$�3�ZF/B�DTGB�H��ƕ%�)6U0r�$���f(hm��*q���&����H�bɑ*;]�8�@�-�b�	 :��H�j�F��և�����P�M0���imm3�mDf�d�n�pV1ran	�MyL�V��\e�B���΀�y�"��`�̎��B�*��i��v����U݂�v�y͝VJ�N�-�ﹿs�`Kt=K%�$#�"Rh��ߑ� �	
����Uc˃
��ut<�7R���K�,$�(��,I����*��lB=�U!`[7��,D�x{_]����NQV("�0W-�A�s�se�ګ���1G��2��|��>m
�\(%lX$A��+�1���#V�Ƞ)�n�BHaܳ v��^y9X���z�Ԥ�*��t�n��@F�!�ʯ�BEF����g�-ђ��c&�����Sh�{8�&:Ai�uT~� ���ra�0$� �Ie�tF��a_��)�x�" �J�5��c	zc&�!�����ZX*d�,�!ؒ	Be\J�u�_���o@�g3d�$�I����D�s�{��75ᳳ��Fv�SrrBR�̂�������c �vW<���$�5�E�6�f�Ɂ1A/�Da0"�l�(�Y�Z��KϐBu��Q).AFWB�݂R��F�r�	,�-O!'��)/n�g�
��1�Wļ�8G���#�RDy�8��A�Ɓߎ&�A'c��c�s��p3æ���r��L�;�)]��l��I&+S�Sc]m�EXR�G�:ݑ�clM�[r;�:�$$(T��P�0<f1�ť������%R�{�.q`ģ�(��k��И�֖�p��')&�6�j+)ǋG~�eY%D��k����l9�R5�7*�f���J�w��:	���mM����2�<m���*.{Y��J�$,a�$oq�?��O�R�_���U��c��T0�R�R1�M��koj�lp�W�B��p�\8&�Ǜ�K���3�9ҳ֓m�����r��T �3a���9��*��&��dC� �����/99�6{��b��d*P�1�zc �=��9'}�a'@�5�g��ѬP�1���xOF�1��p��J���~,`L(_����lQ�����!�aM
��h�޸�������B1Bq����$�2s�FI3�*���	q"�-B�oz=Bv*�G��'&�f���쯍hF��u�2D�$#H�J�P+�D�k�Pc(��^�� �L����5b�"�����B"ȧ�5_9���1Ǌ[(�:���� �"�ݙ�	"q ���<��vB��[��\6��o u��q�{�_r/n����*
�%�t��bd��޵NbB��c�S��e�ޑR��tn%[g����� x)��r��H ���&rI( �݋*�����$k�&�.����γG ���X]��&h6f.�RwBkpP^��C1����ʰ�uk! ���1��HJ�)����+�"�/+PH:���N!��LgWbFm����D(Q �3bN1���C����a]`!���	@���|
-W�'=�x)	vUUo�鈪!T#��7�б�$m�E �05�n$�>v�>��Ŭ0Bg3@0p���������x�I�� vS��FCo�m��B��']4�,�<��;�
��Z&B� ��{H��$���gi�M�$�B��2��֍W��0RTt5M�f;��$���l�0&�������TH� ���Z����.2��\E�7"Am�ݐ1m�1 p�"T1�r��=i�c�]y�d!2�TNvc��g���B��ְôuxL�p7YD���\�c*�w3*�2��)B����>#����&C
Sc�f�A�g��m���e���`�3��47�S�V0d@�H67&%X��4���FSK��إ,�yU5%A��*���&�����l�l�ؽ��ɵ�8��f���B:���\�/k�=�We`Ĝ�;�H4|/�^����-� -���vn;�ĐAx�V*�P��B��7?��1����KPwL���^�Â`Aތ����sK�|y���)%_\�JC��w@��)r��P��H)���/
w4��PH@`M��M�B�f0�4�{SSL&P�2P���m	(P&b�9w�|q�/��G���n
o��"*.�ӏ�3��p��XFe]h&"_z;u�n��F��c��Ow���R P���c��{s*� !�{�pJ���<*�%m#$�vJԆev<.*�����yq�����C�H�f�se�N��=Z�L{.�rP�#Y$�g��A70��0���Q�S��k��A��nY��x������:�� �҈�[ ��iX��]������:�A�&�WF�	�$!��Fj���w�B��yj:3��BL�B�]��!�_�&o3@�Q�<�}�D�^E�b�Y)C@
@����!��ŧdJ�B�!D��]� �"�d�dd�Z��7M|���!�Lb8��F�zo=�gt�1}�\B�.2�V��������Ȥ�D���FkaHL��Rh�R�`l���pqa�Ǔ#c�`���DD��(�4,�u����6���|:IB�-&�,d�]�y�6�90K�U|��A�%K�$B�s��&�r�d�S��*HÚ4��5@Wz���PX�nV�r�D���A�D��!�� ٕ$!Cs �hojC%�3�����jJ%��{A�M�=�߲n`m�dm$�a�8��f�^�|s`��sB��p��B��oQI"@��D�E��F��6X���*�R6�Uc��Υ�«@��f�AIP�^U
Q�!�a�f�\��Sj(X�y0Sj�"�*}�>|c��ʐVuV�W��Ղ�8ƀ�rOr��2_�����0�9�3��\�5{kTm��;���:ܱV�B��tN��07�X	ʈ�3��9I�Z�s1%�ZՀ���n҈Q�0��#@��A6�K�t�����mP��^#"Գ��A=O|�)�-Nbq �1��X�����`��@y�N�6��$!�R<�����@����� b&��&�B�Ě� ()
��b�\/x�� �R
{F��	�!!�UD���żf\n�"�0�aT@�7tX����x�3�b� ��d�nP��"�b�v�͓a#j�L<8��ݥhlLH�@����tyH��n��+�\X�����@0.n*l�g߼�S���n����%}�&���۲��qD%��DEΌ(kè��B#%P%.G�wx?e#ֲ��=ϳ%��A[#�\v8���RI �I%�"�*[;+0�����z�#�L"Y�lAP������
An���ɮ��@E�^;�\��c�c�`�y�B���D$c��CEv3�:�0 �T;��z;�s�t���׮�e�F����7���340A{��#�+�|� .R�0H�*H"�^���R7�q~S�R)ݐ�"�13�T��I�
F4�B"�h�"�|����H1�7I&�v��R��$'y�d�QH�0B.*]Rͭ�_�^�\d�Kg**p�f*Ό�7GN�H�(`��4-lڐY�&0�إP @B�g��s��n>�"�H%pJ�8k����&��N�S�t�/�)	�q,y��5�)Ő�dR��+-�Z=B��E����2D"X�5�f���/�0Px��(b�$5IGm���$�XT�)�G��� ѩ���{f�8Y����w�$��@�ڪ�4�|8�&�X �9]�clȀs�{���B���"%"wBEF�]bE��Y*T�d�2��.nd�X��(�PQ8M�X�'P����I�).7"��m��zN�y0O��"�! aR,:%م�I^�R�H
,S�;sCغ�Q	�2A"�	2�&��0D�DĂ	M��@MP�TB�L8A�d	`"+b��l`M�%�^�s�:���NH3ޝXh(:@��'�(�[��X����eE �J�H�{/gӉB[�ڍ�D�(�L ��\�ᙏBYDZ��p0�%��!��M�EѴ�.D���|%�L�0��l�AƧ����Z�F�!j�V��Q	��@��!�n���o#8!���$�NeKU8y�%v�CdB�!	� �)]F� 6��X�A$ T����TB�BC�AP�@��
ɉ��n�^� \�r���`�!&
c�.IdD
H�I�b�T$	�%J
�f)	���9��BU@��L��Dȵ�#�c�U	�v����4�P����کSŔ)r)	V� {����-�el�A�UE�"�(�PwH赛�[�Z`�X0pA�/0�*�u�[�ǻ������$`�\!b��*�!~R]�/��|�4fq{��B@*��(Sw)�	�R���
D	$$�#%�e4"1�ڊ��[�A���G#��@����Np*�D�l�A���:�0�59[��R0 ���(HK.ꪑ�Кh�7��q"�@80��!z��`�ܬ*$b
���ږ3$�]Z�9@�J��Bvv`�H��+$�qF�ɰ�"��b���H,�!�L$�`��Aid?�K�"��V`!D$l,`-�#��y�&��$�>�#�e�=�����bL�K (�Qa2�hy<q2���1X�E�V��"R
�%6$���أ">^���8��d�5I�
�e�jA!;��q;Jb��ܝȔ�A�A	�wB�a���Z40$��6M�	�Pv�#FU`�K�*����#V6l��3�R�!�(��0�?r���L��d���K`�����C�t����X=��#|,8��J�Eb�"���4x��*�2(/�ܒX!4��k��Z�D�3�M���3EP�#�������$-b���
��0@J!H;^��fCJ�1S��Vᗮ���	J ��{ �^mt�ѦT)!T&��i0���q/T�L�N�.`Ȥ"��AEh�勃=N��]��Y�1b�.
��]P����"��K�^��t��+��*�4��#�d��T6Y���HƗk��Q;b�lڮ;�귋�3J)�(�:��ڑ$W�Br��Q��:0|=Ԣ�Y��igK>�A�22$�~��pûȋU�QvF�+*<Y��t����b�8$��X�H���e
�WQ|(dekY�2-V�$*�9vSRº�+����k��UP+��vمU�Evt*E#	��I�=*a�A��q;Vz���B�QWx�R��F��."�b:�m�E+EP��
��8P��2��
�F��
A� �蠝"��!P�yw#�n�[R��de�N(6�ʖAʈ��U
`����ek�P�EF&G&7��]��+����,t
�MQ:Vn颹�o�۰�h�f�9�FC�舄����M�˗��bV�,%ȕN���E	�,�WEc4��$��Qa��ݑu��˔K�J%ܵ�=�T�����:IQێ�H�UQ���B��=h!�&JXV�Cs�9x�@�c�����.�(�omє#�4][~����%�ww�Kz���a��\8܆�)G�X�V@�#��XOFʡ�1����8����K��S9���`���XKWP�F˾v�o)�d�H��(`�T�fdae����#m�(Y��YyEY&��ᱫ	lCͧ��e�T��C;F1%F��$Ϣ����=�<�ْh�Qr���`��V-�8����ܸ(�H�"��*8�Z�1�q��#��K��L:0Wfe�:K*�#D���م�ED%.�\�� �K�U�V�L0ڌ&������!�1�#�"�VJ-Ѧ�$ȥň)VD@��U�X`/>C*v3v���Se��)�֒E�M8	�bL��ccV��)c��4�q��-$S���k�A�6�7�3�AĆ ���l��e+J�	X�*�tbQPP���#Dj({�9e�GY&0�U捂!8߾*b��T�qk���R/3,	l-4�Uw%���T�=�w�#�A�Iڟ�g�8��AeO�X��gC��(��	(�k��uԎ�Y���t���dh�sd�鄶�%(mk��(kB���*6�u\l�􏬕�a��7l2$��*��j�orQR���HϽ��,Q��+Vj�0�$d�D1=J���T���7Y3\�R�D�y�d�&�@UV̝�&,1G���f:����Պ��~�Y{ ��:����������a~��#i��Z�"3B�b
9��^�p��V���N�+�j���G�JQ�F��*�0�4�.J���rf�: ��B�Ēd�D5��i�o'�U���H��#˺��1cQ�+�š�!bl	�m�J�ý�<�����XVS�־*�Dr�Xv�Y_��u��mZ}��U�Y���veeb#�8�p;���\N;e��Τ�Ǆ��j[��m5�in��!���Ԩ��ڊ�|g?S�J[�ne�ɱB7P�FYE��k%�6��,�D�p��e)1�ײD�B9:k��J���,��`Lc��h����b��`������\'�5s�y���6A�coqM��%�f%Bc��!�������~ǅd����YStD.�U\�p�%���	�] �vV!.�����̳�茳��[�Pqb�B�Q�d�4V	F�t�ߙJ��t5�&�֨��2D�#u���sQ�G�m��ޅ�B!3��R)����H�:Z4�Y�8�/���TFyk��U^$9Ce\,��QI��y���J�U��DB,$x�j�I�-L�Ir�ff%
�yޕB(�Z�1C�b�u!o��֩7�Cv�ބ�bm�
����'#ځF� �aoSi6Y�GM9f�D{�/D5�(��yͯ��E�3@���U��`�&M�'<�n�9�[�9�'�Z!�[�w��bL$�Kp��r���\�$H|&��"���[}��b(�9��H�i�Lazr�1Ld((�
آ��YY��n\H"�8�#�ؽ�
�Ϣ�u2@�^�D�U�I�=A�+3�gl쨗9��0�S �A,�W@���\�4������'�!9�b�&�Xw�;��K��sm�#�� @�r�V8���^�ׇ�����֍Ù
��eB�69��=�A�BL��gB�F�ʯ?$Y���/�<ʅ$F) &L�26W~��o&��Ix>zY�Ȣ�����ˋY&�.)�a�������e}�
��
�"����2!��L���; 1a`g23Zŭf# mRA"�?&u�%�s��Y2d<H�A\-ݭA�{���#w7)&H���'�6
���S�K����es�F11�����*s~c�f�̠a�x��ǡ9�=q���~�?V(m����3>�B�͒%� ��u�)�BĦ�|Α}霄��$$U���m��!8ز0`I^��m߁���x̆1.��ͅdg��M���;mE�R,)�aX���H.����H+�����xH��%�d��<�F:N�˹��W�eY��%�$��Lt����H��dʕ)��^t��("xh�I8����w��L�X��$m�i��i2�U5d'G����8+^��J졒�r��]K~e�l:D[���!�7��y0�R��Ε�Β�9�����@��Y�W7���1�,�z$"��C���l�cS�B�M�K�-r��*���~B�Z݊G��d��
E�fI�*r3Z�d� {���qlZ]2�<o��ّ�a��FQ���D�v�n�T����)DqR��`MP(� ˞�������7#Y�����1���4v:�Z��b%[�S�d�E�Ʉ︳�3��agE2(F`̘���#��<k��9��h�P6��J�0����p��I��p��\����V�.̒��EH��D�2ҡ�#L�R��+��۾ħ��3���i">�CchXZ�N�xDVWPR��wD�EX��@��Y�29R�X��:m���V��T@�j�H�m��^-�.�s�*��TIV���#��ٷә����R��U\l�!��E�K�)��hD�|�!�A\��"4����FsK�8�c��<.V� �J���h��Nѿqv�*�f� e��e����3��u9	�aM qQ��	)�Y�0Fj-+�*)D"�J+X{��Ľ�v����P��e�.��SC�i�藸�i������nʜ�٥|���C Y�@��.7�'Qy>�y?�\@���/���Z��7[�Ǭ�w{l2cH��y��@Q9��`ז�������Ք-�a�����!R#�P6�){��X�@����(��akY�k�Y¿h�\^��H��7<r��`�·u��Ae�[{��K�NB" �����T�e4�%K�m��x	�|��-���I�eL1�����~�%{�Z��R$�D�.U��[搐Q*ܒO�
:l��FA0$���B]BD���:2���A�p��Cf�ҨґW�c��p�"�0�����\ i(��kw��{��T�/��#b#<F"I�Y�rx���$�D�=��& ��}$�"���q����ub�[IՕ��P1��&�P�&!hh���Y�AK��x��R�v�
xT&��ˮ��dWY�M3%�NJ��Y��ټ�:��uL�
�!�0Ad���L@wbU��	�h[�Á2������M�����đ��g���Df$	�n`�����ͯ2�I� '#V�ڦ���"���j�A�<����L\��YBYr�$IFwK'AH�Q�<6���1����EC"m���\���8��_� �T^��m�G]>O+�}	���7�#B$w���Mi�4�a{��R�+��ds�eX�b��aV��e�_i!�lK�"���a���*	�T��awJ���$�6��	y�2�;��R)�h�"{DLs-E3z�m��ʬ�dю2X����f�v�r2a�35^Ϩi�r��������۷�웘�]���܉oӠP���5i}��k�i��Bsaq�g�3x;��7*��x������:��2W��|�$�����b��-x㊾E�S�� �:D�ERNdAU<j8ňRSck��f�����r��N�͓�F�@����FUB��N���� |iRu���%!l�䜢	�['�Q�5�!į$�/"L��b�
ܧI?>�����`dB@��h��7;�j�)�Е��H�zQ%y	<A~{cf�N�Ǎ�ln�%�m��c2�*!C�Ç�$��+�X���B�Z�Ul���P��`dѳ�'gJwK�$E��$�""IPXs�Z��;��0A޸�U�0���p�{Gl�1<�,��)�ZE�b�L	vf�]��;�n�X���c��0/�ٲ��3�ߊp5�am��w�P�F��l��8��{RY�d����C�9��=�m|V֝�A��TC�E{�q�<����[0|�kW��*�@Y�;���������3���PXP�!eA��Z�"�W���

X��6�R'���ף���x�8L����؈���)7)
W_"}���
���}4:~��o��Kf\ �����;���+���Xj�	�$eoa���HW��$J�iL�"%B�C<Q��w��0���A*#D�$	gc���c@�֪�F�1X�*�|.(���0DM��h%F���[��ak�!�7"�A#6�S�6zE�=�v�	� �Bm�;5�sn���p1h�G�&�	�����c����ý�j��\�@��D̓��{V����� "���q�-��7�T#ĵ��J�)(X��>�{m��晆��nR��DB�n-�q��!`���sw ���A�H2n�_���Ftۻ�CQ+��DR� �*!����I�����;��@W��:C@��B�n۶-�Y~	%p-x1�La:T�dm��&
D�"�H!H�	@�7��,0���)�^u$�4�XQR�A$�IJ(	(k�ԣ�j��ƫ�(`�U
(�R��Z����{�}$�+p.L�W=�����N��v`�f��Ёt<��Ȭ"��'q�P����U�^0].�[��ML7���Ղ9@A@j���80��'�V���'B�
J�ݠ�Q%}�cC֤u�J��#	^'��&�Bl��{_H�9�g1R�Hk�8�5q�Tk �8\�N�3"`B�j�+i(�d~�v� b�T�B	0%��0��u%j��aGI� wD!�c�K�Je��Ƅ�4P�: �L�D�%H�"�8�ִS����Z�<�m�Hme�w�����0��Brʱ��!2�%�V�b(��,��7۶�Պh�i (���\��/On��1`��p�H\����L�6��,4���hAR�F#kE��J�(����:�J�;4jH���SA �G��.A.V�J҇U� � %Tږ����h�����*���CCܨկ:!��DĮ]�:�;����X��S8Qy$�[��\���B.�p&7�]�����*"I�(�����;�/ߒ�K�� ���Z#J�O�I��B��/g�!�(`���[�28W��)Z�K�d �CC5a����ByG	�PuX�ra�A�"�z�yE����5�DҀ�(a��*�]��Ņ�ޔrک`�@$*���f\wJU�ÇB�����#G����sB��4(�(T�\_.�4U�K��W�pa�� � r�� J���{HE�dnEu�*	�J�����S]�6$��Y�Da����cP������U�5�C{l] ��m��ڈ�dӍ��k��HV
JʺX�
���KmB$Q��hݶX�!5J���b" qH��>�$9���H�!�0[99�2�#boj�
Y��f-��jh
?�� �;x��*�������(F�]&-�i1z��piPR$�@,C�QT� ��g
<�2(H��s �cI#L&�yHZM9(
B��	�	��6nkCc�-d��"�'��/��2cg�*3[('�Yb!mcBT��'9�f�0����0�x�g�)�M1�1!^�����jȓ�(A$�0D^j�6����甄�D�iSh�Dl3)$��D���C�ԑ�q;���"*\��J�	��5
��t��!�5�Ē	�Ŷ��h����Ųv�P$�T��"�&�"y(a
O%fA.D.V��9H �}OAP3tC�ET�X���nE�M �
�5Q�̂@�O�Y؄EB��s~��FDm���=�.6�)(U&`&Qu�:@���]zބx"�A@`L+_�ƣ~da��P�6�:חg���7x��}���&�"(tfˁ��|�B���l���R�Wl#�:`Q��4q#�� VţtIM�#����):
���H��b��*aٯ=�5��1����f��9@�qW$(@Bi�����`I� �\�d���#F�$ D�S	h(&SP�P&Gц�9=TbhIb�d�h�`�K�a���"SE������d�L�U	]�63Eq*~�ݲ�`�rS��Z�H�pQr�wW�W �)B��`�
��B�~�1�,�K��z0R���Af2� N�Ss+�{�5ԡ��P��,�S93U��L�P$���mw ��&sMKBJ�m�(��Zҍ:AM*��2ks��WU�X���WX����$/�%�WX@���Z�B;�D�è�����X�[g[�5uB�:M"9r��VE��<�.A�)��~p�ƒ��T�@�v�>ͣ�8�m����qu�*T�F
��pX0k�rqV�88 �2b��)�}��hP�ZeW�XXeE��n,�O��D?a�4	d�^�d���L�.�D����e`}��� o �����#JD���5���w0� ScPHx�$-zA�5�܌�1۫<vH���2J�24�BQ�o�Sg�	h����{+k��t�rVՅ���l
(m��	@����o# �,�4X3�����n�%P��P�ʠ!p�)Y��bDJ�(�IN
z�43Zr�h��DP{�n/"��ڵ��@�atɻA �9\�!s�yΫ����TEcsÁ��AS���d�{��)@A(P�re4�(�]����;" �ĕdj�F}��6J����Cx\�	���lv"Ȃd�I"G:-�F�eU�'�(`��$��ӤYV��#c�.��B"	�,Q_�m�5���!rf���z��_JL���u^L�-h$b���(�R�SI"�6�nd���[3Q����sK���j@$l��@�@�
(H�3z�p\�N����g990��`���xZ�K"L�,m�I��{|F��R�S�o��#�V�		BJ�~���L��H0L���
w��\��id���ͧE:!H�$m}�_j#��O���I�jB��D�l�!��a��6P��.��Cs���@=an�A{F��NE��0�kvIL�'+��A d�Z���XDE�ۻ*�6A���r7��A4I!n
"Dd!yh��XZ��'�Ff�(�dP�t��G��禀jYI�F��(���y��r6ŋ�٢n^H��T#�e �9@(W"�
�U�`�߳7i-.���	����`t��ҩ�(Fn��K�d���j��F 0q�3�AB��f���f�U�!AB��B��p�g��:.�$�UB]o�`F&�L�D@�Ef�.����VXUTm�W���`���;W�@�3v+W�����̓i Y�E�]`�H|�U7E^���Cd�JSÆ��E�V�E�t@U$'\�t�*�Jܪ�B�,�t[+EO�T2l	{D� �mRE�ڣJ�)�.�+��Ft���'
�3�V�AKUȱ�.�W��D�����h�3eG���1[��(���/] �͔�-z��DK���f�F�Q�����UP��I����9�f,��h���
� K�dgʫp��ك9��ϝ���s* �@�
� B�*(H
*L.mi�R��n��#�:���`���ۖt�딨0� )" h�DWn�7`�(CQ]��2�*�*B�J�� � ���w��r+*	賐��A�Tݗ=�� �Q�D��<�� ��7���G^7�����`�#7_nm|%@d}���+��� �;�!ǀ�c
�T�aP�!(�,�@�(�$�H�@(D({+�C��Q?8���E���2��"J��S�D�{]\��������V�c��p97�8!RP �A=���r
�D�� � 7�� &I �Av�
���K����0 ja�,��	���z"��^��t@t_����f�v�C�uG��|,�o����{��~W�>�������@
/*|�U���L���7U��;pBH��|��ݗ��������π_��8��'���>���ijx�W�OHa�z| 'P�����(����`��� �/K#Ġ)�,Xz@ǰ���>�Q�����ܭ?�1�|�DUMX T߁Cǉ��dX�4&�2UЮ\�dmGJ\�nZ��Ơ��A0�3��b:8
�4�M08#��d�&H�;�QAEt�g���`����*� w̻-��\i`̍U�!m� /��=�ia�f%�H��*(���`�M�n9pFV��z
��[-� :$��쮆����`*�c�ESUMa�[�  �C�5ɭE�q�N.K��$��"I�S�s}j��=$�ĝի��I��I;p��w\�܈��/�@�<��VEHĄY��INF^��w�2��<9�"�X%���AQa 'A�IB�dIK ���"D��_Z�뻣���׹��.뭵dWR�zOb�'����5$R�ՙ���k����G�h�	�h�-1Q�����1��py9ٮ���0f?�8�aw-3g9��Y.�ƻ�٦1�l��u��9~rN�sWI���6��u�g_]��oF��7c:�d<��%%8�i�\�h܍4��ad؀� 	�K �(ܰHIMګ���A&D� ��`�zݮ^��Y�M� E�1�ÇH4s�7�7 !��@�@�e�@�	�T�]q
(A��#)�'78t�ːvi��F�5�"��,�V>�C��%�8d'�'⬟��3�̂��5�^�ɉ
 Z�b1�C��}�=���CR�?7�x�����?'L~�F��#�>�Gu��Ck��r�.��L��� YRJ<(\t�CB��� K��@^���@@S����l�h
��l���M�.-�&kQTD1���èg���<=4�Hp��|RY��N��3�}��7Qی�n�"
;�
!�sf,�#B��dg]uTCST7x�p{��Xuw Q⇛5c�{�X�$���g*�a�PF�@QÏN��H�1`1`��� R9��8��!\Um��	�/�\�&���v�� )i�8CT����"H�P)B
��͙�ɭI��JkE ��E�7$:�*rwM�!��$ÜV =L�9C�u��0���5Up ��:i�?}��x�� �(�'�!>N�l��ʢ/������`�Hq1\�&za��~d+����#��!,�
�	8��ˡ�E�}|c��2�T�9G�J?#�~0j�B4��vh���g�s��:X�k������E%T�����d�;��ֿ5ŕP_��P��]=��8���O���&����\(��L�G�'߆ S���vN����>9������F����P��[�����
�-�vM��~��E{��z�f?�{�"���'��D=A���?G]ϵ��I^@
[G����4����Y�)�yL�+���(���F��-����d2> �/��@�?��|�������w�������g����>�%�������������@�a.�J��!	)����t<D\��3��P��1LIh>` �-�vl1��@�o�p���X� X
(�'	�P|�'�gD�w� M@�3�4u"J�i�)]��PP�HJ0�����&BT�lCx!���<��i:���5�s�nz�t!�����=�G�I�#�d-!���C0��}+��"�A �S�|H�p�C�)C
a  Z���w�7�:[��܀��D<8���S���NyG��~��(1�ܨ�  U����ju�
(9��8ǡ���~L�UD~� �`6�T��k� $��t�̻�D(AB �-'�wݶ���Ψ �x�#�:�ۂ��&�v jm썧Պ9���� ߕ��u��'���|����̠��A�( �fXQ�̎5NV����Ҋ�
dv ����J{��O��7QGUM�P{��_�����=p*���AE�C�v�� �Щښ���5	RM��|
'd ܇�{���t���1���8�6�E h��j ���w@U�p;ܠ�w�N�]D{5 t����l�'�r���N��CE���ӫ��ǟ����Hꤽ�:��X" ��[��@xM��]<���91�z�\k�+����C�܁Χmх��ѡ�!�,�KÑɪ'	��BA�=�t�!
���<G4t�Ӏ�,p x�r��9@)��G$@�?�\¦��Ȁr^_Zc���k��-aC�\�����
{l(��B�<�?�����8�:aCi��:ƀx�SxT�#� ��0�A�I�r�uM�q;7�N��v��gt�6wl� ِ����@!\9���*�AWu(`�\$!��$�]>H
cj*(:���qP���r�;�*���v�A��5/��Oe�'�7�)��:�=P�E���8D���B�xuC�^ ���tN��P�:��@9D�P��H��.�]�ɨb%HIu]���C t�Ԩ9C��9=���{��p1k�xo�J�r:8���5���L�
(��A�:WD0(D��0��H���hCpC�W����Pv��"�� *�q/�C �*�u�CA�����=�cn7ͻ��3��3t^�U�����?��D��Y r@��.��p�#N{��'�@E�(s��7�FE]^Z��*����!�x�|������4	��<b.���h��vq�-x ��X;p���va�c���>gI�r�Rt���h(a7�w��E8b�����0������h'\h� ��9��'�>'�o��+��dD_�z��<A��O<�S��z�wF鏞��� �����pe������C �����'|=U}ޘ�_��4�<� �~t�����׈|f��#�d?Y���H�2��I�?s��uOsW�Q�=WQ��CX�ސ���E�G��U�9V�J}��쀦�����c���F>��$n_j~�c'��E�
.n����@���߿Q�=���_K������z���{����_K�}#{�~~���<��~����,������^s��������G��;W�a���&��C���G%���V2;Q��?�\3���>�Y�����?�a����K�җ���N~����>������|O�7ٙ?�2�}���;���J�[����\w����\ �����Uz�~���9;�s��H?��11�A�_���~�暧�>���%OY ���b~6�������d���?X�����=�&� R ����'�_��ǭ�}W�7���'��'K澃��w?��<�t�"E�?�x�����&/�@SG�a������!(QS``�)�l�Y��_���Xɜg3�9O.�u����	��|�(�k(B����=��M5���{�Ᏹ_���&�C��ϰX��A�����U��OY�y���A~���Ïf�)������x@�߼_	��$p>6?�-/�C�>"e�?����̟*���Uyp���Ĩ!H��?Z$��9���>��EN ;��vJ��k� �u5�s�W���  ���v~��}��;���M<���$��޵=7U���?;���t'� LO�?���������0$����_����H����(������9�ӧ��r����������O����·�"/�WZxx^��}��ڠ�� ~������3�\��$k��L
%������No�]2�hTW
�|������A����!�dnnK ��eA|^��Yb�y꯴P�r�̛V�غ&M_���9��M,8(����Fa`�X�ᚉ�&��.i�0a9���)�����OIq4�;6�ú 4+=-1bn�K1��>1�/����z�׬�t݇v���z=Giݶ���"~߹�bnϋ�C��ǉ(��tO�	:a�M!�;M�C�$>�=P���PU�^�-��> ����^Gf����p�����5�e;1��R������
���Hoeh@�?E%�e|9ڡ��SL/�����ETet��a�	9�DbH��PwYT4 �U���Z �s�S��@�)"��(��"@(@�(@�U�TiVA$YT�`�HVP!AR��q*���!�� ��
�2� �+(���@$�$ �H�$(*�)�
0!
��
@0) )Ȥ ~W�B��r�e �3��g�Z�����˕Χ��uηweӶ����]����7�$�C���v��O�{�4�/7�g�r����w2�,�%�buf�v����n����ݛ���|�7i�O�����}���!�|���� 0��� ��D���3�%�7�Y<�9���4�W��qZ�,����[�ϐ	��u���n;g뤺:���GA��t9�OiS��L������1��M��.�Cc*�ժn����ɽ��
E]���$��3�y�Qݽq�"�던f#�޳jᎪol#q��h�oFEd��ӧA�7WI�;��5�f�ݖ틼��ʒ#
�H��*��
,�B� ʰ*B	 a RL��J�ԧ������N/*V���|$���eF��eub���iV�.���D����o��^����2���zVd,T���6x�^LFF^q��e��2�IZ��,įiF+��bQJ���=�8��mG��Gt�ҽ��:�,�Ť�eg��c(���E��V�G!첓�Lg4�-9�/w��{%��[�>�j��c|�ƹ�H��&��%Y�o�b%��])t��Uĩ�{�mV��\�%[M �  b � ��?�<.�����cP}��xN&�%�TW5��c):ҷ���\D�4��ҵv��W�r��v�m�jTo������d�[�带�E2؍�5"&|�
�gm����I��k�em��n�:��zCG|c{���N9���+�q�P[6�Olͣi�w�M��Z��2��]��4e���l��x�z�mSl��fV��kD�F%�m�i��b�������z�x���lo��)֭�mG�[d�4E���<<�8����j���l �q��}S5~6�˰s�N0ɭ���īK��z�Q[.��V�$�Riݵ����qx�f���n�|�jJ�n1�\�cZ�VJg9⯗�b l�ޟ��u�Q���i�]w^[��ۯ�	S�3��G\��;l�n�g��۝��)Y2ǿf�A�ĵN-�b7��ｨ��_tΣL�'�������������-���Ӟ��=Z]�vƮӾ�w���ݸ�<v�cn���T����Z���ۻ��g�Y%M�E��.���B��Z�E��N7�}�^1�7�n5����=O{�ɿ"}G}m���j����/yq�P�$���fX��]{�)�#����Q��HS�U���m֖��؝yx�:�~�L�H�Ws�҂Ϙ��-����l?h���!���);�켛���¼^�ݻ��N���۳w	�i��|�z���؋s�}��Ξ3��_�#�*;�U}vM��O�i�q��[��ޚfUz�n�������x<^[wJ����F���m�ڝ�f�dK�(��WC|�M�"��b��r�ߦ�0Ƕ��6�Yӕ����c�ET�U%PTP�I B�����G:��JW�!,��O����h��ߡ���|x���KcR�݅�_��,e����Yg��=��V�8�|x����iGԷk{T���Ii^����J*:�튵���{-�W�z�3l�Nd��j�bS�ל���%��/�O�/~<��N�U��wM
��>9�jt���٦���oh�c�S�i�Ta8����)d�~/���s��Q�FT�}���۴�56��>#��=��������m�c�����y��Kl>�:�����T9��ZI�-���l���^���[�,���:��n�v���{5�Q���N[�;7��K(�M7���y�j�#�ڸ��}?��?��J�{�x��gJ�=�κ���U����س�z�}�����s�y�}�qЖyU^��N6Ǟ޳�l�8�h9�{����W2����c��*P���Q��=��:��T��q^OT�g��X�Z�{���+�z��~�+�]V�����'o^���_f~�=;p��+MF+ko�q��n{�wϢ�&�)��x�v�q��s��z��ꬃ�o-��V�����V���� � 0�0��V���,b�����B�� H��"�
0"��"�0	Ȥ*�>��y:�7k��x�o�v����{F�T������_G����A��ۏn���?�:zW����W�ԧ>&�״[��y_��K�o���|b�Q�%�P�_Y���W�Lg=xIG��}>����}_�.;}qx�|��ן~���������ﯘ뷻�|r�^�~����<s/C^-oa�9�{<~3��¾3��{�ԣ�ywK�k�œ��}| {�ij���ٽ��]�l=�w��������O��R�Cf�éǉ$�u�O	��'�=��~)`�K�����k>�Rt��}L����T����Z�"��~:���\8��{�q�K�S���S�0=�m����|x����~{��ߞW�]�ߎ17�~;��r���|5'O�{���j�����.�ǜ���~����on���t���{�{��-�p����W���Ki����n~y�k�)O�n'-v��M��7׉��u��%O�=�x|y�>=_��o�t�J\ys�s|��w�����.'�}�?R����^��������g(���4c�J����z�Ez����Q��UŘy4mR�I
y��a4��Rm�p�U AG`S�|��߿��x���=�]���l�^7�w��s�!��ʶ�׽p)߮���  !�}k�q/+������!�������4��y�Ai{#�ymuǑ_�7	�5|��1���F8K�jFs�A��������($M�Q�.)�C��J�(��G�o��ʬ���J�[%�۵O<q��_x����~%�|{��Kj�R�"S$ ț4ı�����Q�<��*��pVt_Q��m��S��������O��k�oѯϞ��{}�G�a��,���F�t�l-�S����m��f8ZGd�R�&�Ea��4 ���PXU����L��0��iA-S��aF��s�_��e���Ծ9�f_>|��㯤���}g��n;w���s��/o�_���\Ξ�2���{g�/\p?>,�j&Y
L.lN9ͦ�c	Ϟ��2�$��**�â:7�aqs��)旑���H ��	�$`A�!`@�n��9"�D�BE<qp���!M�%�MV�^A�*2�,A>>�����ޣ��/�q>Q�������w�<x����������8�R#L���P;����[�Z��*�l��A1�BH�z� ����INц\�KX��I�J1
��Y)�WT�ILdB�� ��q�)M�J����r9u ��f�I"A��	�`�U��Y���C�i�&]�d�4�e�`X� �$(b$�|DXˤh����h��̇�;j�s�.Pb\����֗���,K�̳�j~7D��J�珘����}�߉7���ﷷǖ�v�[�hB �  !ϸ�?�������ͳ�,~7߷�i��4��oo��2�����JJ����۩/�x P
�>��I:���M�7��
�apN�"!&U24�2*��SG��"��@��g�<0��F@9���Q��
 (�p�T�#�x��O�Rq[���tj�P�D��;.�,�:%�Q-��O���T�U��l��X��@YI�����i!���pC��h�m!m%�T�J#�38��8#�������$qǶ�����}C��Vf"碈_	<�ɴ)H��= W��U*�B�,�s���s�*��3����	��d���zva�!\�B�:kJ�I.&ʍ�rI�81�gLb�th�^�U9��:eq\4�1uG�VbEUp$*���op&qE�!����"�
D �	;�LQ�S,�(�aL�[R
 ��4!#�H�R�jl<�1wU����$z�а	A�۳�h���o������#�������K[�~5����c8�?N�����}�O��#��D���I��Ѫǒ^�S�(�H(؋��hy𒪈2s�Ș$Ŏu؆@����]$��j4�h�	9X���IabaZ����Uf��Lm�b%��d/���
�J?D�#��9��(��B%��
J�C�z-ĳ��Y���$�E�yN',Ba��L�C���%�K[�l�Kq�_=c�������i���v��`Y�nh#��(��3�% t���+p=N�8�*ǝ�Q�5�Uh�&,"�h^>7dA�Y�[#B���3�,bH2�-����2p�Rc	�Ē�4��Ɖ��Y�cf@Ǌs�}�}8��z������.�[��H����~����~7�ӽ�T��o�����蠬����KIU�@`��g?�G!W�|����p�Rh�����J��$�����t��1��)� �8�
��fO%$<���Ԧ�g&cDвY�(����фU:f%!Gŕ�R(1a��IE;
q��e�S�
�l�%>x�:̠���Zl��'��d1�Y���G���b@I" ���-�\���E2
JM(j��B��4����M=T��9%RC4�4�Y��mg�x]ԗ�	��2$ ���ԣoD��T�&��%'+�F���N&�眼��GY5��$�PL��b�P�SK�1�l����掝0AC䀃c�dY���xўPiM���ig��Yi��J��+�}��i��;My�;*��,U^ZSƕ�4'��(U�6��
/4L�B4�%P͚��?eL�C��Γaj@}4����(:�. 44(����ay�d�Q��"�	X�#CRf.�	��"(ӣ�Q2��ü+���B˚f�B�l����ha�0u�l�#A��pK1�+&0�-L�Dea�n��-H�"��*�
DI�4�Q��� �Y���R�hH�d��h�݆J$b�,t5 ��c�Z�2��8f$�E`q�~D�5 �B4�a$Ř4�j�D��q.�d�<�Ui��Q!�@�0cp�{����х��d����@�����X�\*��5�,V�t�ƔZ��W� b0�ĢT��*Y��3/�x$i�Rx��<HdT����a�G4�ai4 �[S�(MZ�T��1z�)d�t���e(.&gf�Ȍz��,CnF>rp(�$eo�JH
�l[2C0���#V2p��B7�{h��0Ӗ �p���]8�d�,9�H��GM�]��=D@�I�B�=U��Cd��:�ej�b��zI�4k�G���r$�q�Q���89)���o����iߪz�_��s�?V��_�@C� ! "��¤�
�"J��(ʄ �����@ >� >�@� }>��}+T������M��`ڔ��O��u8��h���mpG	�h��h	I�Pf��������Y�8R��f����u�kh[�CJ��iB���\lQ`��T����^8Q���qB�
�9BO<�,zg�J�
�&�Y+hYn�(��so�aU��v����103E����J�c�.ڮH�+�b�6\M�&��i2�u���믩�-�@��,���]���D��~���"�l4-e�l�2��u�Ÿx#��.��H���ID"��	KY{�J��2��,a�J;�uiRm�ݰ��5F,�"��3�L�Jh�DT��H�q�K���E�U��C���$|P]N���@8��#=��& �S�銉�^H��Pf;�����s�*G�(zѢ��90˾����C"�p;�*�q"^do~��Ȧ�&KY�cPF�Da⸶t��1��4,��;2)ak�m���ˊ���@�jh�	%�I�b���~�p<z�����a%��t�J�����0A!�)���)��!�@ijTP>�d2
�e<do�,� A*-�,���FO*�6: :�l���P�R�5\��%lTM�^�7���E ������#�Jr4��:�g�E.�L2r&������!H�Y]�J:��5��]��VI�����*�L��P�����G�I��i��ZK6
��-6�a`Љ%�H)H�
��1�(�}e�@���
68�6묙2୚qY��dy	�5`��b38TFȍ�V���F)�j���Q50������_�d�uW�)C�S��m���J��+
H����DZ�Iۀ� ]�D��dU0p\z�5�`�&�(`B�f��]��ARB.!ν�T���!�mx�le�_<��cT��`�g ^�~hN�f���/�9Y���<z��4gbu�`hyX�=�+�Oؾ�ڸZ�'L�t�D���}0���\�Hj�&�
�%�D�ͥc>�`��Ve�C�^&�����ٛ���)��9�&M� э
s��u6�n���(��̠�B��zDA_O�>��?�=콟��~c�z����c�|�����N۲�{�v|��s��<��S���u��#GWٹ��������[��/�Ѓ7�����X� ��)'������R��?� ���aVU%amPB�t��,�x2�S�M5�s��!T���6�EYi'�(�4��A�j_��'ɇ���i�y�(��rD���%�2CJY�_ 9��*��J�2��Q#iB�#�Lfl�|� ¬Bǯ�Ől@`�Lq<S�^�,,�@<��|s�X�P�P\��O�܇t� ӟ�"~��IS��!�e#���A&�Y̺L�H
H����̪�6�$�p�A�#��K<-	Y��8Dr�n���K�䋆4 � ���Lg ���0P� r��#&.���xÊA�f�!�&0��TS��!p����T�CnH�!�#")MDFW����!褳�Oa�,8�y���ـ��4oZ���ѕ�-���!C(Ц��s�@��*��&�a!Y%����3�k,�b 4M+�d�l�@e�L�Ŝ�^"�&:��LGDXL�'L��tQ�hȥԛA�QB�e�-�M��d����I���MhE#�Df̌5��C�QD�D3� ��pjH�h1JU�_t�!e��Y�:�;�&�$H�b�m�9ߢ-�2��)��p�b2ЮC!G2�t��Y@�JJ�6��K�W&j��k���imL��!6S�H�|��|ܤt�MHb`�Ԑ �k	dƃ$���J��μ����2��
.
`�������~ ��ž��(K�0Fk@��R��I�R��N1 4�IE���
B�dS@v(4ƍ��K�2��	�FR���uhK�&c���N��¥t�ٖ��*�Q^8P�~���9�͵��D�IL�=+28}(�	���� /i���ڎ��Z�$��9��vy��&��!p5���5�( 2"�0�\�9�(��w�{LfI�,��-hE6�k-�J5�־��������F��kd�u�ℨ��4�������[��UP�m0���jjW)&����@fB�MT����*IP����o��7	�p��\XၰAP��v$?)�g\s�Y�G�S(P`��9�!nF�=�UL�����@�Zr�mM녖鵂�f3UL��¬�].[.��M�h,�V��Aaqc#��JgG����g�ZA ����Rm�S�F���:�c���N����ať���9�Wm�N9 �4� }>�U:c<�O��FGYN���0���2Br�Uէ�RK'a����)�[P�k���er���0���p;�Vh��v�hsL39%�.�0�W�sI�	Cx��@C��ɤf�gY%i�x�e\�ӆEN�\CS �c!���v`,��)%iK�M/R����v���"�A�\�J��(��܀i-�y�����!��aJ0]I�=�6�T��#�"s���-6�KWa�M;���)���.sU�����&M���N.pՋ���Y8�L��`��ﵑ������ː�+Kp�dQas��B�&X� ���y�~�C����i�#\�?��k5B �x��vО�!-�7���(i�}M^ĳ�=�o���d�RP�=&�?	b��J0)���{�Z���L�4NuU:�U�VN�RI&2W{75xf�=X%�QH�ؿ�_�=Ay$�/^D�N�)a �$���Z�ߢH�Z��a+=8ii�,8����K��"�#YSU��Ա���J�t�"`�;[�\a�:=o�P?��V���LjU��x��)ö�eC�U��c�:0���Sl�B(l����Y��gl�6�M�ǖ��z�L�~�Xx��v@�t�;O��)�Wc�kx�AYb��TJ�x
�.Ah�)8��ݗ�dTK0�0%�OL�7=���r�N��r��ycL�����X+F��k+��%����T<�E�y���WZ�&	ZJ�%ۡ�A�TʉFi�a̶���eM����M4Ť��:o��W�R�{^ZVI`�]�ɇ����\��ј'd�#U�Y�a�Ճu-����H�-wc�7'�o���X6F�Y�Z�Ja��]�bI d�&��h�Ƈ<�u<�G�QuG���y5 dy�ۊfY�^q�Ŕlv���V!��-mhh��� p����}Q[��hKgsDX��i�.���3i&�o̸!�:�Ѻ�^�2�Ҫ���Sr�Ȳd'v,�`���O�-����^�n*%�'f�pn��&�c�����Pb�ua��{'�y�^��>�g�sc�v�´ !�4��|(�3H��%�I��p괚cyӁ�C*ߒD�aU�,�U�Dg���6j�hj%Au104����øӬ��Lf�q��w�Y!�X����*���t��:V�/�NG2��(2�{߬���L�@�!����j���Z:235�^��Қ�6�%|�sC���A�S9�+��r��X��]���IZ�DZ�c��W3��u.�G_�r��g#�9��Q������_����7��f	��3�Xڵr���nQ[��-�
�DW�J�   �F��@(U�B���C3��4ŌF1\�EF6��'w�����Ow��U�X� *@T��<ł�"�`BR5S��m�@��ݔ�כ(�]�����r��ޑ�.c�zm��Z�5�6@�V�Th�V��۔��1���(�h6�Z�'����ߤ��|?G�����yoQ��;�ޛ�����כ����������ө���f0DQ��f�ceH�ґ�iB)5�U�b�kQmREh���$El&-�eZT)�*JD��)P�D�����(����V-R(*
PJ�m[i,VѰT�Z�$a��
X�h�!D��ZV�J� hU(@)iD�i D� ZQP�T
���T�B��)�R�)T(��)
P��R��)�ThP�PH	F!J%A�������W�L��"�������_���ǳ�|�������/�����?��������7��>��~?��O��ދ��_����w���G��hB�1JR�@ vgh�����V��cL,�����3(d�@&Q�&@��)�A�L�%$�e(�d��1*	 )�P�B�a��0�EP(LLE&&T�e!$���
�`�$�� �"#S""CIJl�(��c)3#)E!���FŊ$�1&h�R�R�1$,�Dd���B!��M#������O������·���|���ߖ(���Q�������]������{o�}����yR"?��'�~��z�z?[���N��S��{��w����=w'w�y^w��������{�	oG-�$�ʕ�94�3��S��R��5���mQ��fj(����[:j�w����Mȳh�Dg��� �l��2���JC�u�Ul'T���D��Þ�'K�n�0a���f�1���G�mhw�/�BNq��"�~4���Rp��V8,�D<o�*�+�1/�&I`���tl|'���Re��4��%�@���KU����#d���ۥ��E6�ul�XyҊ��S�,��"ALdm���K���7jY}6bD4��1�k��M��zy�V�9���g�U�8���q��{�ܒ��dZ�%t@����f�<�N\'jy'�V��2�\e3%wJ�;�,a�����iG ��nY'� hf�q/�v_�T5I�Z�~������*;�>+�!�:Nפ�����0q�ͷ;�Ge�� ����O��`���A��,�����a��3�J!�)����E����g�������G8��G{2Z�EwV�bfַ�����y�C��``1�4�\Zԇ�m�LE)HJ��n�2�y%�f����d(B�AؔD��`�d����<L1�YJ���Bw$J@" ���$�έ2j��hc!g�z�f�P�	a���'��)�g8����=8]��#{����P!��8��NPMU��3p���MsA�U%/��ڵ���U'�c{�(�S2F4D졃W������ܬl��*9�;����@���{&��:�����&+lHڌrǉ��m�wR�a��� �x�m��q���ż�V"8@2�6�>h��tM����0N}#%&d�Xak(��g(��0�?)��y�E5�ɥǰ�!�jd��& iƂ�A|Ҏ���m�n�'$��:3/K+�:�v���lB(�4m�#o)�ަ��ؑe���mܔ�a���G�RO�16�R*s�q����nՑ�f�Z�hk����aC�q:}v&*��ل0�}��=ۋ�P˦x�����r" rLcQ#���dMH`�!�wDwP�z�I����PL޻eU�_��BT}>���P� xx3U�Ї�%��I��,��}���>3�I�2<����˦�jk9a5\���-X�ʭ�d��sj��H�^��}{E��$"jƥ��)hW��iǬ`Q��(|ݤ�;JƱ]�,zo�s\xv�ȚZe���s��Z��yW�) g���s;��v�5������J�!D��p-�F�WE�*����u"��Xg�a,�
��0
�Úb҄�<'n�Ed��S�?OC��ݭ�b��5u��8j(��3Suk�a�iJ�a�2�AyD>��ܲ��.=7�z����\\ο�x.�u���w�F�N�:�?��r���H���>s�{�Y���a1�F�F���i!����@��wY�b�d 3+��&�\،�@� 4�0Ѷ�.`ݓrS0�� H
&� m� _'
 �d �TG0 !�TMaA@�EJPR�ZT��V�Q��jKQQf����V01�C~R�l���:I���%;����Cdl�%܁�yT1"�SY�2R&��@8��g�UA2)Zk���e5�׾�p;�������������������������������������W��m�U� `E�;�   w�L    �              
�     ��           � �            "      o  ��`                jQ�;� V���y`1�N     � AB�    �(   �mI@  E�� (P@AH�     �� -§      0  �`     !�
 nX      rP(�ܻ�  <      2IE�    7      � �z�
     �h�                                                            	��      `     z 8��E��� "�@P @                       @  (H @       (    P           ϐ  !�l �-1:,@ � * h     �   H    s�|di@  4 @} )**� �@   �      k�C ) �   �     UO�       (��ɦ��0h)��M4�(�i�4$�i��FOS��)����zjm&�(&�4�MzPi� !4$Й522hj��&�H�S�I�S�P 2 d��SA�   �4  �   ��A��h)S)e��h�A��L��dC��aL�@�A�4h4hi�� 4i���MF@Ѡ����)T���!�L &&�da4�`#0 	�� &&&F	��2d�т0`A�  	=RRQQ��m@ڀj   �� 4 @ ��h    �  44�    hH � 4i��&	����i馓� ɡ�6�~L����� ���m4�l<�0L	��)�S�'����!��z L��h�ԙXd�c�J��d���og�xN�e�GBA|�{~>B^�Z�%]b�0�˯�abԾ�@��� -�N�#$se���`

e@4U^� 0����sW��*�gCP42m�@B"�����/�����3ѡ��(1���Bp��2XAU  @��9AW����L�Ù݆q@�� (J:"�z0�e%�d���*���ː��V��b��U"QpB0*����/D�T/]ۿ,{o�}�KW��:�L  QD@�8���Q�� 1Dh��[E!!'�h%R �[J�AC1m��V�i��%nl��iѰ'�,]E�S�� (� �@b�5�T�C��W<� ��`8<8���"&�xS2%YK3"�  ��(6������U��l' n	Vս�W���C�����q30fST�$�HD����,4�DDOn� TM	ޫKX��o-)s84 ŉ���� �)jRhP���S�f1$o4� �L�K"0�B��Ě7e@4`�	_� ��e�
R-�_�m�-g��"��B��M,A����6PZs
�hv��Ƒh4f�r��@�(���.Jh�B��He�4l��T,�s�Z�;8O�ed(��1T���k�F���E�a7��_�8P�$��` �F�9�6\<�_����FS�l?Y@ִO%�f@X ���Ѯ���c�X�ˁH>��M��YB��Tn�/r�(�ڀ4]�g�7�R+�n��=�ŗ���a����j�lv�
v)��G'��+Za�pl�9Dچp��@�tr,�Z�1)����r�eTZ����Tb,P6��`@��^W�Z'4L��2�m!'����\c�j���Ljv��]2Z2�ZPX�f�Ul�	�HG��b����lYe%
�z�g%��p�я����B:��u�g�]��0�2<��On�p|��h�S���=kv�֚�q���*��B&Vm8��N�Dg��&(
�>P:**6>���U*�B�} �V
�6�M���#n��×��j8z�.F��������}o����$�>Zā��״eUI9T��<4}�p�̻.�Nհ���j�`U
���oO2�=�X��=�?aĨwn!
m��;1�_S�jd���J�~�����G+�͞����)t7s`�4����"�yN��5j)�D�{MV�,��]3�ڌ�j��p���B/E!h;ޕZKeZ. �7��������&00"t#ezF�!I��W �B�l)0Ė5�6�/h��)cxF���"����8��70��Lm�QhXũY�N���/i��������"����+�Ea`���`��3���m�Qs��B1S�#��#Ϳ�����r��Tj�Y��� �iҊ��z�4U4����h�����@3�(,7햗&sf?�5��TI�YB�<i ���x����,�m�t��"��#���;Q�
 P�U�B"@*��ep�[MHͱ����yW�/���[�*]��N/e�qT,��pX�"�A$z�������?ϥ3,C�mEEN[��	��ZKiK~��7��\�L˩W�䗗9q,�m�]+��7��>>+������\�.��\�7{�	I���ĺ�n�ȗt�=:�z�qA�׽�YW���緓����j��V�͋���5�nQ��6�ɵ�Q�i9_-��ޣ�
3I�z�O��EQ 3��|�BLL�۲R9��մ��v���ޓ��K�|T���@�	b�yIKYO�`����	��e�p`��e��}i�d	b��%'�3Yj6�Yj�Ͷڶm̬q43�m3&��k�6�6�q0Y)"�Z�i���΅@J��iTa#V�Hd%�kjP%+/�KF�����v6�M�lR�V'��5<�
��m�5K(a���F%���D�tl��`�*���Y���f>�����mW�b�*Ņ�� g��V/�_[TKFz�/@Q����  r$D �@dv�s?����FvtRI�$�I$H@��-��u�x��Ȉ7�:P}�M!"���E*��&R�@
�"� @ 1A���@B!�vX�<N������Q�HBE�U*���PU+AR�`�H�@ ��P" �E* $"�(O/�f�l�L @���<* @������"	�@�i��̃����  }���O�����������:�����|����g�>Ls�o�b�s�|���ߔ'9������q���]'��t����/%��������o�"��V>�� .C|w��/���~x!�=Ie��h��������ҿ���?"=�%|#?0���$���.���z���9����H  R`  ����=!x��+�N�m�P�E0�0�@�{��n����a0;�����O��0�D�"��+�m�HV��N��˵��e7@�����/S��~�R(�ħ��_�o�=tp�Ӽ�k�H�����&;Ϻ�0�1��l�E�Ed�q��;@� @�<�"Fkl��Rs �um����{���p?�_�|c�۷Ө 'h)��?���� a�'B���0�Y�d@���@=B4__��l�)-@D &w�/�;�x?������	��Ixq��)K>�x^&��ϒ���4ď��e���<\���暢���}0���_�{}� @��ጉ��1 	��o�+�56�c��v��� �/H���u��k�5l�1wiv�N@�%��Ī'>�ߐ���$F�����@"'��	Z�g�~et �1� 	x}�6����D���4#� �"�Eun���/�M��1���7D�$�������f�S4���" #Mc�5��?���a   B  &��q��w���������ݛ�y�g��B��ӭ�ߒ� �ol�"	�[�!�Y��d ����X @���v�b=���;�����le ��_9�% ��{�^W_5����oL������Ӟ` O����&��L��L��"DE���Y����cFz�d^�E�n��Bna����^WP��3�
�48� ��ݳ�v��  1�S�/nW�Ƌ�K�gR0WD"��������'���,u�|~���� 	2� ���[���43�����^�d��@� �3�0>~�1~���7�����F� 	h��c��h�hۅa���"͙Y� �6�u��oшiC�*�~� " O��1M�W����6ϟ} %$1]��7��]$�+���A��Z�W���:/q�|0�Ǘ�D@�|FXa�?�N��m_g_%p @�y��%��<��z����P�/���R��Nڝ� $��+6���]XY�(j����>��>7@'�v��~�.vo���D@���b.�߁��k\{x�֏Ѳ  "3�y+5�v=O����r�[���t*�  $�mx������s���6}<U�ߗ�1x�ڊ�x��� D	A����zɈ�a�6�" )��{N�/���x�޺w�""I��P�gxC�Gf�� W������]s��xa��� ��0����q���" �.��o������Rk�� H<L��}��3���D}�	Z�B�6�;���cG�^Ӷ�?K���f�w>'�ڜH�:������˩K64�+�q��x�&�\l�9Ѵtӏ��==�� #�V�<�ţ�o�Ԫ" @��=��B�~2��� ��"�z�P�81/DQJX�y|h�֩�U�p��Y��1d����e26��cײy�%�<��Rs8I�Fc�W�h�ļ�LCkz�
���]B5�j'�����2�<(��D��=��_�ʌ�>�JzG���[ۻ������":[8�����aX�j��M6�e	72n:	��L5���=�����0�>I9�,RDUu��R!�>>�3�,��A#Y﷭�z�	�Ϩ6��'���"m���ӏTXIJHH1��m��@��ҁ&11jMpT�["-�V2'�k�>���K�����mF)�[}}$� �o��C�5#+�cz�z�O��n˭Q��x��_s�g�c�0�$H@�$��]֙���h���x%�@�Q�u�� /Fty���� �|�(HR�^-  ��"(xX�!��IX�ڕ��&"B!�<��IIHJ�y�f;�v��!ů�>$:�rB1"I8�Ы��/c�\7�·����ʊ�g��%Zz����Y��keY_�m-�]+��Ve�ciaXx"��u�]8HL@&�ǈ��q�.����(��!V���i��0E�E�JI�N�ܖ��IR2���5�1h�uՄ��y+wY���h�<����R�1iG�|C����DŽl�Ac6�u��[x����Y�,JBkv5���=tӌ2����a!^Pǝ ���a��lZ3Ɛ����*'�����u���V*LN��+S̄�@����a�
1��B�OD��(�,��̛sRQ1��Q"x��޲�$S¾=�	�n�"k��ho
�T��D�H� B#�R>�̇���#5M4��(�/Zg��Y�2�]�n $��$X�gkBkl �Hb`,�Z� !�d���4�l��@+�6��,Vp�� D�ŗӳ���Q@�ǭRsk�k��!��k�����v���9�N���e:�>R|w��a>:�1 9S��im�e���	I��R�X� זeՖ#��st����Q"�X��+�0B}����0���RS�Z�u��	Bc���Ԑ9Rhx姱a%�V$T�F�Oq{/��K�Vh�	ǌ��s�޷�{�Ͼ'��cG��|{��VZB���wY|�]�8tP&=`�!	��v�5��s��ī�>;�::Z\�1u��YW�>}YС�=ƳX����jK(J� V�	�6�B�	H��=W,z�r��Cֳ֗��Հ��U��-o�W�[�_m�s���,��=��[6��R[OR�)��J�M�Ig;#�K�v�x����7NY��a��&o7�Ҙ�8� ��d���j�T����q8�Ϯ^|��&!
LH�>�DJ�F$RqLH;Qx��&#l�B��RKI���I�Rsp�բ�LRXF�Xl�yį�o=^�� ��^;�z�X�}ǒ�X�'m`a����
[{�zᬋ#�Ix�n����Y��1�`���k D���si3��l;��ϩ՝�qLC2R�絤D�ӡ��]`DB�}�<*R}P��lnMb�ϙ�dDA'-��Rll󔙈�����MDz��aT:�����t���_u,���,�;q1�ǉLY��W�6�y{Y�a&S�]�S��ab��z$�
F'�f)��fWktH&�T��=O���T�-x�`�i��������<zC�׬�<�O�1V%��cC�)�2��[�Pf�:�b2�LR���aa0��@��hq�R0<B��T�8k9�ij$O2�U�LvS�r�v�9e"vq���l��L9W�hFve0IN�ɡ#=m��z�x��!�r���ĶpB��]a�F��"�#��6�ԫ	ɛ� �Hov�=�>�Zݶ�:s,)@Ic���0�|�9�x����,R���BT�gr�&̽��]X�pfg�N��z�W�wJNuCu���ψW��m���*zY��q��%�Y�Y�A�H[q �#Qd���Z����# �R�]x�F>	�s;q O=�!��t����#�+)�X�=p����;y.�M���d�Px��ezg�D�<�O᳗���.��x���D鐒�iS��&�`c�%�[_{�A�V��/I7Y�{��kܑ�ڜ�8rR�l�8l��ސCL��%��I$�t�VvSx�zE��4GЈ(� �V��"J�� 6p �F�����O��a����e��т�ba�Q���P��aA#Ye;�����n�(�^���G�gmx;@ N�_p�S�f�.���/u�|��,��e0�Ǹ�́1))�#a6fO>c�- ĉ��c�T��Hf��-%8���<R��>�� ��k1�ޝ8z��j��Ǿ�}Ou�
}m�)��4.<0�Rɷ\�쇃xV��$��<)		lyƊHD@H�ll'F�[��w3�
Lq'��/�@�u�~�)zzY���P�.;N��<x\��X��BL�b�1HT$o>�%S�P�!ʉ�x!�V��ex,$Oil���P`�q�6tg�W����<z��-q���s��g�A1o�$.���fg6b`��a�U$n�wLC��$+�F���/��Ԭ>�8�!0$!՗������z�Sʮ��&H��x=�h_i|x����ǐ	B�J����ԉk��2-R�x�uԋl{���-Q�퉲�����\�ѧ�bSrfJG�y��6 �y𑇺�륥��`D��8���N"5��g��;4��Dd �bK��ǻp�˶�D�M�`M�̳IeV"�8������ke�����3�D��}��f��i�K�XF��c8׬��FT�I�J������)��igm�He�
>ac��	OXJ�ao�!`1)/�=*$kq�7��t�,�ɫ� �6�LbN봌�}`(Ґ��3�|h��~�P���ܾ��bDJD�mP�Ϭ`XGЀBRF�яoj��b"��P!��8��z�sB��8����F�� ���mL�:[δ�� #(u��
�uqՠ���&y��$���5���IO=��	/�S1������s���I��|I�����\!��b��V���1&,Xߝz_x�R�'��R��>VE�g�?���w���O�bo�}���o����/��n�������[������w����?�I'��[�6����������g���f)7#�$��1_�H�)C�d������h�s����Kh��?�Ҡ��QD^���k�4��5������G3ͳ��xo�����G�����w��������G9�/�3O��C�����_r?q����t���򨯽��E���<�`?}�����߷����W?�����;�w�E����yz���Y��[���������`|/�歟������#_���w�{�\������2b|��ڌ�O�rIy���z���n~��\}����'������������O������S���?��R�O���d~�����������i���� _�=϶�?������zN�T��!����C�ď���3�G�>gĀ�J(��HV_�}s?���V?���֐=%Z勜�ڸ�	e@�+U	2$���x�&��R�-���|�y�u�O���]�x��o��[~�j����`B @ ��!"�$C����#��b��0M�}9��B�T/w���!��$����<s��Ї��5�l����5C�(��Z!��pW۵�tm�P �4_u�U; ��0�+���[lOA��E���=Ǟ}�ǧ6�\R�m����tcДxa*�'>�ć,`Sݻ�'��Z���ؾ|���`��JARG��v���a*��A��L��1
�}4�]�Ew�K�7�l-e $ݥ���j����,��9|a!�a5�U�p�"���|�k�!-�B�_nhQL<���-\S^i 2ѕ ��
���'r(���]ڷ��)�'��da !�|y�[��[���tu�-�=��4���6,OV��8���.qKZT�ؾ�M�Sٌ�^��P`�8aA�<�GS��U!'�(�RI��0K|��R��M�H�|�_���!9���a)��ǂHsI��olPW4�D�H#�-.��[/��2�ԍ����b��NնM����2o7lRXׇ-��u�Y�"��@����6G�6�"��`�3d�𒗭�J��B�������L�0N�o	���ڗܶ�Txff�aĵL���.�FŔ�@<x&����XY��!a� E����[{��i�J��2�neV5�X���mb�*O�'W�Y|@*1�B5�����f�RU'c3�-�@��=䊚2ؤ����Z�����'�
p����l	��I�NZ�!�v�d�y�,Ys��\�N�D�>�\��^�n{;�ק��6��� 1��Ya`⬻����6z��`^]��>�9�u{'�ʲZ0��1�=����'1 ���E�'�f$���4woP�}��&*Z��z$L_6�:ٶ�u�J��e�B�v3	�VPa�<�q�QH�/��lK*�U�o�  b�o���}�F�c�E������X��;F� ڒXNR��l��ta+����a	��B�oWYjQ"�Y����#gϩ�CԠJH�9���R�|@���V���ńy��	A�lV�{��C2"�X�YO$	*�ȭ �֓:�R�%:��1�(X� ]�ۏx,����i��=Ů)H�z�O $d"!� o�l�c�1{�%r[�	V����Ȑ�z�к^,=eRB��,�a1�bi*+���2Ȭ���ql`!:��2����-Z+AzW�:��,��^��)ھ.��x�����R�}Y��S�	Owm4}z�љ�F������_z[��)Y�A���}Idz�Q��Q�E#B0�YaY������h�%���+| �D��.mAR��Kt�*ȱ,c �m��d NY�}(/��YI1�g�T�B��Y�� �s0O 
.%8����5����fԘ�!s�Z[l
��� n�ǲ؊C��!e�qJ��a'-XQC����� C�f͎���a���gY������1�Yu�HG���
���`�<DB�����F_V>��ل'BՑ�3jb�`/��	Ik��i%0me	D����aI_4xp�(��ů�^c5L���:���R� H�Ϟ}�*���X�H���Y�h.mcI�����1���Px��s��Rb�/��YN$��QH��{��x"c����-@a>'�|��BR#�c���!����^]d"�q��כ�Qk�����L� k�K]U@fRP"{�z�U��h'��@�^"d�F�3�XLS���}M��P�������	s��q5�g� H�o��K
BQ<�Ҷ����X>B!�����>�Ј֊��a%�1�d�^��"z\�J��nZ�@� �1�㬖�D��H��BJ[H�mJ�Q�bT|�z�[e���m�z�a���vW����zc�*x�[�1i6t�Of"@V3ǅ��01F]o:_R!�c����vq�Z��{��]���P<y'YT���cE�'_bK/��x<���wN�q�]7�_h�cK9��<u��b��;���8	����ŖJq7=��+�B�U}kH�ZE�c<B:�en�*��+�}b�P^,����|*x8���LFVcs:��^RZ@�s�v�P	y�&p[��b���
��0� $'uj��Q ا3%sƳ־�� "�X������W� +X�����O	D"� M{y& @�ARsl��k����w�,�)-��C�Xm�m	Η�!
D���)� �-e�n� tm�9�Z�z���9ĠC�dD#��!u�a"ua X|ud�2�������Ǻ�fTG��%$!�}�Y*��MZ�Nu�!Zx�x|ί�/����g/�cY�����keu}(�[,�Fu����ǔ�lР��u��XVM}ۋ{�u��]}�'G�;�J�i8��9,���X��+����H��|KS���zhHIH��c*�](�=�Xb�ᄧ��P�T�Ω !3-Jx�D�&��8�RKNi|������!oi�g����È�Q<B(N`��QJp�i:�a����hN���b�)Om��6����c��6|
��T��c� ��+-r�Jz�)9�ι�X��2��
�IlR'�$9�ne�����<���� I$ � Hkk5�鮶PY�}LN�"�D�σ{�q%1�+����m��<g^�����P���B+��l(@��cCG��:P�&Wq/.��3'�flI(E��X�q.:�Y�[5��"�����M9��傢V�e�IH���m�YlS`;mBN(x�V��)5j��^�-�w/	�@y�t���r�R�� ������q��n�����T�̲��!è�s��j�j&z,�_R[`�
J!"A�-x����oi�R�$�8���!	LX@����u��HI�3���	��|�
ƾ������b��wY|�_ZG��D����#`!��M�nn\�*�՘OϢKlb0��e��B��X��mo�b�OB�`+�/�K�%�0��}��N79�^F�B<�V�h�Mf��T ��5�}��ǡ��ς��S�HT-���C[���ih��� �Ĉ��|ф����pT�<��>�t����-aR �� �d�T	����{�9��w�y�h��&��jռ��s��{0��ľ<�Q�WĈ����ϴ@m����ؾ���q55���uB��<��݅���������me�����e:�ւ$s#.HޮO/����̪���)��-1펽3��gP���$���x�&;��gkɭ�馃.�� �HVR�ф	/�!���-��@�G.ݩ��f�m��P�F�"b��1a�ɺ��X�֞+�Hx�%|��ֶ��1,�G�͸�"����؄֧ފ	蔆e 0/
�k�,߷�C�{��$��O(�TDR�E�D�	E+@4`��#h �(��</n�5����h��|�ߟ��?oQ;�����7o���˰����ɖ�ì�������+�?��E�7�?z-]��k���8Y�5����{  � �� �� ����#�U>�߽Z�Rw칭,��őC��ɋ[��kTYS�H�g��;���
W���<Q�!��-앥��vN_"_�݀�lgT�f���_b����)�[a>�hNɇ���[���Ѓ���~E@��L� F�c ���Z��!�$�s�_����o����m�H���{�ۉb��2/��x/;�d�a?QLf��j��rX;�S�neWK;���Z�V�w+�`w�;��c)АI?Ҋ�YAd�&>�9\����B�����.�ɕ2PHU�;�L�,���&�:�#��*�ʡ<�1)��]�|Í���f�r�CJ�'�P&�^&	O!c���9!
�D��b�غD�Y��zU�Q�Qd�<�<eqd�J]%$�����/!�r�N�>��)�iF�5�	J'?��i^ů$\��I�=h�{eq9�ҕ� t�X�+� ���Fs�{f��b�)��b,|�-e�d@p_5�EE��I��({)*�8&�4���S3˒Ѳ�
�д3�-τ��R������o>o��+�+MN+��Ք�D1<���-�������Hի,�|���̃N`5�se�S��%$�
�F�)I��TU��`���������&5&��K�RB�.p؋*���q0���G1)d���0<�i�׫f���5�7�u���C{�pSSa�<����y!<s'B!W�y��C�F.����~�KD�u�l�eĐKEb@P밁�{�哱����&�*V���aa9KU��/ &d����[y�$\i�v'�g��ISf�:X��aI�������P5�K=���fl�.mF����F�
gW�E��jR6��4w�H��wrR�s�f/�6�S��8��k��OИ�P;��,as6��kir�
�7Y�Z/;W0��Ô%��n�cU���_��2 �o-H{�ͬr�R(L.��P���Mk3�V�c��4��$�#����c�^�wjOT	t)j��mDݻ�ۛŤ��Ղ���I2"�N�Qr��H����!Y3�[�ZyȾ��SHjk۝2�΅��E��6�X�V2��B����uN�I�w���]J W�Ո�l7^��,cP�1Y�ߨ�#��P�٦��hV�A���D�\�'{���ڊK~p�i��a��3�3!�{4�]�U;�`��Ez��s0Zk�!wd��cEP�%�����O4P�ʗaS�끗P(j��c��h��`I�W�ս�����sq�)�p6�g���=9f	��{C�'�v��5�x�TU���lz�ɖ�{��:nY�1ɪ���&�l�b�}��&ʬ(��5Q���*(I����u��uuos�˘�%%X�49S�$�)D�<�v�0�4!a�fƄ�:<Cz:�hP�Y?Q�aH�è�$wuT5�X*�k�O��j	�ƞ�gRI�#�E�8����:�
�P�U)�^렃��B M�2���ߤ;n����b���7Z�ކƷ��~��&�s����c�vEO%iG��Q�B,�#`��aPU)RB�b�"~.��t]���އ��o�����>^��?C�����_�4��CW_����l�{{������q#�#�����1����fO�)� �:��	`��/�~L���ߺ��"?�γ����2M>���Hli��^���6dI��C[(�-�O�z��`p`�	��|�&6?���46�qV��e����I4~�	�41.Q����
��+5u���5-��m�	��0��m�^��2�br�B:q׫W�0��԰y�r��w��L8������+P�)�䈟�
�H�[���x�K�zaI�j%<��eNi�Y
9Ȍ� ������<�d]��n����J
k+$¶��>��9��}{_0J$o��8�=6�L#�������OX�l���:J�vAI�u(�鏌�B������)R�����	�xK��x�I�O*�
�u��m� &M�N�74n�=8M _s�27���t�!d ���(aL����{���r���os�#�p�"k�|�OG�
�O=��z�ᯕM�1W��/�����dX�ǌUq�K*���\���D"��[��j�P�P�P���V!��&.Sly��7��l����3/7đa )�q����6�D�-��qxV�r��*��f)�=Q��7���E� R�6�=�Hk�EҠG��VwE��vE."y�y��yF�Lc�(�f�:�G��II�����F/]]\��]��E�Ȝ?��*�ɽ�Ϛ�Y��v�#2D2�d��J��{K���C�/y��^ f�J�Dq��A����dQ褡&�ّ��G�b�ZRY?w2��k䜲�CVR��1!����XS�z���_�XYZ6�W-�������^�hV��?(#�A=DY&#���� Ph8��:�z}�,Id��kT��k�D�e$Ҕ&�#B�b�9�n-�!	���5#<I0�6y���mR��&r%�7��5�:so���𩊠�O4�%&-!�d9���i�I���*��cy�A0��E�y�������4��cë��	��E��L�}0"�&�L���T�FX Rt�l��۫4��O��$�Y��a]����H!&�2>#S43��с̇Pu;��2��-�@x�-��B��Ul�u���D��o�r��<��{.7[x�����HX1�te�t|S�4��:D��䒫�|����^PI�`�l�!�{�U��n"��6;�x��q4^����uc�T�_��[C��y}Q�輺�?w�p���O�v+_�~�+A���Pæ�v� Ҵ��DfNu~rm�|˺�bC�K2G�HDd�Ht2�R�ԆB�$�����$@`wKEf/^sQ���ʙ�V�DeT�	�-��M��a��2��n錒+W�Gt�i�f�{���'ρk�N���i��&&�E�MsH��+�Z��B³/����Q��fu��:KF�}�sM�c2�.p�ʨ��*���u\O>�>�ŷ��6�ap��玃/�9^��[��S�ѵ���Ed1l�::O����a	�b�R����7��P)#z�>��S�0��xF�G���r�
؍��WgT��p
�D��]Z()��C��:�MuRWf�h�<,H�X�B�1��JP�P�sm��QG8�GV�9�@	�~&\Ao��m׹����J��H׏<-���QQAm��L���w)��ZU,b��'YE��t6/$��j<�J���=2i����<"S�c/,��Pe٧B#�*�P[� �J)����#4�ryi/�8�Ժ���4x���#����$���:����AR֊D��	�0yf:�y S�PihD���F}����q��\�/��cN9)�#6/=�\��G[�C�Ý�"��-v�y�M��O�n+�)��4��&��8F�L�t��Xْ�E���K�ba��Y���	k��Ȩ��Dȱ�]�{��I�v�Z�eV8�U�G���@m@q�9KSu*%��iJUYg�G6��q����bi�B��A{�W��}�>���S�Lr�� ��1Q��@-(V4}�?o=���;s�~�����+(~�����}�*   " QY��S���XR@d E������d�c��jM�����b�����͋lD[�t�ڊ*���&���6��Ѵ����uȣ �,! � �$��"�������w�d@@�*�b�
")�T (-BD$D�a�&��(B�n�h�!l*	r`� �X) pwE�(,Jp��ve�* ����SJq�TH�	T/	Tj27@�R,�"2"���NN (��S�v$-�R����
u�Z/!�@@Z�&�`�Z.��A �0� ���Ŵ��xr\h�,6 
���*�� �� (�dQӳt�1�DQ�%BE�9�b�-Pm2�h2 ��� ��jM��`٣�SPD��MTu�*:�dRØ�p��+"���T�M)�$TQԕj*
��#�"� +�\#�V��4�� /�̀���&��D�Ԡ�Qu�#�Sj��h�հ������:a�����6� ),GiKdlL������� !@V���KZ�P5bZԂ���(�j"(�QA�WP���[E�Tb����XdT$$@U�A$PQ���!�#P�"��"�B��,�5�-�H��UVƋj��Um�E�k5y�Vܴi�yY�mEdD$�4�Q@h�����*�"���7J �H��1) b�Ѥ��H��(R!QF�`
�� *�ȡD���V!d��0V dE� ��d �$����( *4�DP�ETH{�~W��΀ ���256�,�Z5��;V��,��=J�H@��EYi%B� ��$TD$A1��_l2cD2\�"�V����k��-˕�k��V���Q*�薊�n�������h��PU @Q�� ��B�U�P$@�\ڍm5���7+��^TW�߁�q�I��[�GE�Xś�y=�n=K�͡:6Ox=KG���bx5��E��\P<N��Gӆ��_%W�-�d�	�>^'�2�Bee����k(|�h�����e�o����3m���{u����Uf��l,S[�lq��l�����=P-���Y�h-��O��A'�@���%Fp��z ���*�����<<���	�ng�:m~퉂%���������u��ym�Jx�
&��'���~���eA �Յi�>קs���ݻYX���"�A/���3�6��
u<׮�>�����󾴔_���Ə�$U��e)(��}��p��ɹxIT�*�5�5��!ͪ#�X�����1?�l��W[�i���#1<?4X����A��O���?o��R��O��XiF�wrcDE<p�Ne+��f�z�8��)�[��C>��ϥ_z�@BfZko[*H�JF�Yh��E��x��aD�d�"��E��6�xL0j��M�@��Y� �kC���j��C�Ř�+����!�j3���X�)S�Ѭ�'�j����4�!"s�BK�VR;O��1u�~��}g, q��Pq�O�7��O|}��a�ye�|��0��0� �-<r����0��a~P�$=ݦy"x��H2�S�)8j�c��F%S��n�x$�iH�!�ǋm�~��8g�7ƌ	���"W�B�J%b$Cʰ�VF�5�@	�a�[c��gi�b��[�
V��y۞�inx�sZ��!u^}�,{��P��m��or�j�)"P���<Ml����ug�f�<�K���us�4`Kf�R�������g��u��P$ڒ3���O8�[#�`�lT �fe�"��	-�)�e�k h���~e�~���2�9�=d�X���}��X{�5e$I�zq��<択��a�Y��4=^�Ѥ���x��%=�ʠS�t��g�@&���Yj/�$=	�/����<	�M���Egu��>�ɖ|=>.�s5�j�\�I�YCK�A.|�eG��zĢ$�	����v�̳� 	��ؚ��t�RR���B��z3�� x"��|$:#��ϯN8&z�	]����,H���}� x�V��� �Ǔe��>���	/�Ђ%��䗙eJKU>� P��ݐN[)ap� sIp�|�qb�_c��-��XJ<şY��[%�Z8��b�q-r�
R�ix��Ƕ�����[Z���[��'��_�c��|L{���>l��_����gk/`�:Yمqd�{����P�1�L�8Պ�>RPY�X�����K��!�1�|�9�12�ﴳ����9������:S���#�tuׇ�ɹ�s)�6tX�c���|8�	њq�sFF�����ٰ����z�O�)_0 ���q��;6�*H�z�Ҍgɫ�)�bk}Ko:�Ag�4|@��
�m���>'���I�)�c�}۵�	��4%��_R��9}2��#_ IG[*ʴ
�5��!Ro���`�0��@a1aǜ��Y5�3yw�kK6JN�$H�f�sz��������}(�Vg�hO����v�#�C�5��la�w�:e��Ɵ6�q��k���V	$�@�o���c�H�'Bb^�}_��)a <�u���t�����\�`�a`O��+��<��"B֕�k2�/�V@	Am~�ܳ�/�\�X�!e>��8�|��a�6�Bg"JͲ�`���8e!�	�a�=iO�ڒ}/�ta����_*���"D"�Ǧ'�o����@|��&{���
���	I|z"���I[ǽǰD+[��#����V�h�W�O0��b�͇>z 0�O�+ $�}�_��Q����<����<�i���>ǩ%qu
�,!~��iH(DVN,=���z�'�Z@�����%XQ���ĝP�ƺ}��<��T=��0��0��=�f� ��`sx<��e�e�)ͺҾ|HC�m G	�����׽��� �W��_��:[o���n���( 'Ǭc,
�_����V�6��_�����
�J�`xx��-�&c��Ǵ`T<|u��@u��p��f����v|�{L�XC(�KYHC4��|B��������5�gıc	y���'�z�O��x��e)4��V�a��jL�|n;[⡈=x��wJ�u��V%)��1kD��J�}i�Xy�u��@��,+h{	��;��{�{�㟶�>�}3�c	�7���0y�;�|�X���am����s�l��)+%��0�Sŀ�lo�qK�"�~��r��9Z���aVYݷt��Y>7}i�>�_�J'�B[��`|A_�O�;��t#k�M��n��f��
j��~'�N�Ĥ�%�3m�kXz(����!��H׉(��J!JX�}S��)V�8�$/��$��8��$��$��'�I�~��H�_ow�b�^E˚��/5v��U���^^^Z�K��/*6�wqlZ��ѵͽ�8@KZ��_�K�}�X��T<�������U͋nmnm�� dq!=b�$�D�1 �� �!�P�HH���A`���m��U�U��� B1�O���W��4$�J���p���2�?��sE��>�+��E��70� ��#h�Ф�;���>_���o�ijv8ۂ���E�d�����"(?W|;�e�գ�ju��V�O��
�y���ky֖;j�G�Q��?��d��6��K��������V���o���zΫ+��n��Ȍ;�{ڽS&��� $�������n�B��-A��؁Q�UkS��6�H�FH��T$I�,� ���*5 dP���=��|$��OɨUT��W#�\"=���I{�Y���d&2y�Q4����z�Λ��}����=ʊO���_|��ꂷ.m|���^�0�S/)�� B��$�U�P�c# �"S1j(El���#d��ZaE�\`Z\®���ZT
��}S�|W�\�>Zto5s{]�^}/)C�7��S��"��(���;����&SrFQ3�{or$I��wH�ĻN�8����{W��AcnkU}�V�V�\���.Z+�k�\�K��_�y�:V1{����]^14F�q�$��9������t�]wq���Ѐ���aM�\�y��.�M`��\�I�H�6��W�Dj(Dd�7"Z6�TT�|A��r��,\撟�-XgҒRD���"��	��Q{�����;� BI9�9q��#�9uܔ����nBI�v�-�ݮQnm�<�ʹj�T�) )"�ب�EHa���wW-���y�](�W1�
��ڻݼ��͹w]s����ǻ�Σ�����wn�˝΢RD溍#5��uv��H��Q������<�9�,�k��#b�E��P����I-H%����K1��:� �.WKsk�N���#n�e﮾-�0�]wm���ˈ�o���B���˦�coz�Z��Z�#h�T�dd$?��p]��yݿ���;�?��ҏ����~�>����?������D�L��~P�E������?��_���:�/�%�ʁ�՚������Oأ��`k��Z�e��o��Z>��
�ܰ|���Ke��K���s�rT�A�
�A�I 6�r��oњ�\�j������U��8A�.�e˛��ѹnwq�b�;7#]s�r�u��ɋ�]�t�i���E�=��d;���tE�rQ9�<�I��~�mZ����Z)CH�=_�f�����9���H��V�����v"�����!%?��Ѯ����6%"U��ȭݚ!dG݇)��c^E�~9t�t�7�����m�ɯn����z�-'o�7��|�B�LE�Ժ!�+{x]l������]�H�g��[��k�/���2$��# Ȓ#"���ई0���4��\�=���E�M{�4��ts���6#rv�0�7:�hl|�Fb�������M0kΖ��yni(�#1�&Ѫ-EQZ��Zm�����(�r��:[���m�eݸ�e����"�<"@"H�b63�	�t\���ݸ�78b�]�Q����@��!��>���{�o�/�������=�A�ao���W��>����2'�9�>��_�ц�dG^���nզn��X���jM\{�0���Tg�1��G���T:��B}�eOl6�T�Z��m>gu���z�s�Z�ν5�ڮ�������x��3��n�S�?ߚ�B��*�н=�WGP��3 'F֑)�d����}�\[m�#M�W������Pu�
\6��,�5�j/ �ަ=5醫���ġV���[4��n�%�)����!Z���<BH�2��G4|�m�-�[�=ȵ��ɘ?���`�����?ˀ�f��c2{��
�[�e�/�]�.�̚����-͛���\�=� %N�W(�+V6�\���ڢ頾a�L=l`�IU��C�n�"�������n�l�)T�:6��������٪\ا}�;��޷�ayZ;�Ā�`�rq�X���x �["�1B��Ș^�78�`������Rm��y��@�<V/&Z�ԍ�T�+v�^T��������r�շJ�t��|�Y�U/cȑq�7Ǟ������D�q�};m)r��a%3"���P�\[i���=h��I�E|�ٞ���WI/��%�6�.��yw��I��F�;��&����=�(��G�_(86��n�Zb�W���X�Uc/�J6�<.��(8�'\-$�Z�p����c�|bwe�꿙���+m��>�6�E�.ZjƊH1R�y�W���raj�C��fkc��<mj�׊4���I��,�U��s�_�����!�D�uR��/ų�5�F�8���t����ælg�l1���q,�_�S^4q��%�ö��ʙr��3�"�~)2�IȔ�Fn�9%㽨v�o>��"
�{�uU��C��׋b������;B!`�a�SS��O�8�;�غ@s�Qv�j^ւ*?����ס(�ਣ��-�jmc�R?�A/����WT"�l��͉�2-���\�B�h�I-g�ض��*['c�]N57�|����+*��h��썍��F�	��<O��,�ϾGT�BƤ�G�%?%6�7��J�e	ıY�]{b����*��^��u8˷sg�h�#ǉ<#]i90
Z1J<�ՁN�
���	Wk�Xvֺa�:�xA[�UQku�2;dw�H?�yaSO#�J{o��f�N��+kn�狉U��y"�ٕ� j:7�u�!W0wB�uG��NaU�"q�7#������Ts��Xu�濵�=J�D�����j�s�wwwY�_^�&J���8��`z.(y��9i���p�^��BP]�",�C½��N��>#�Ҏ�N�3 ��b��NF�q�LSS�ΊǞ��͡D�[Ҽ"�慢��g��Y%��4A'qМ�K�|N�ǲH���mcE��z��y��u�,M�,�(]c�o	��D��N�{�U�*��+(�uY��e�D���YZϕ��K#��Uz)(<�J>��V0�ߓYj�� ���f�ж�+�ϰ��zB�E��-g��m�Wrv��>���UO[E4���T�|�wK���G/N���RS�*ߚ|��8���d��~�I*I4�RpD�.%�U��T���K�۾��ʐ�щmRH�+5��2�`��I�85d:��]@�h٫��>�N4�����W�)�u&�$�1�3M�1
#��I�0MB�yP�.����6�d�M�
t�G.��#�,��/[�y�)�*OP���c���P�j)"[$T���s�ʱP��d}赁���֙r��X�ǃ�Dou�'�*cr|���O��w��M}�'����Mb5�c�ɣذ���!�M��ڎ�ڣ��u�j컥�Nߔ��3��7;�>[e�|�T�'7Cb��Eb�n\��ymym_�Z浯Զ��󺻸��W{���Bc˒W��T��I�������b���ws�����2�`{�$�1^�)Bh�2��q��{�F'λ-�E��b�j��ѱ��j�][{^_����V�sG����IAb�`�M/w{������Hh#&�H04�����4X��D��sW,E���ҍZ���Y-�/�x�����];r������[��(H�8�%�"cY7���NF�+�e\Ţ�|W���j)-�r���Y���U�j5T�t�����n�!(Hܺe��!1;���6e{�"D�(��L��Lh��{�o��W��*9��b��Z����1�h�pco�J�|��B��S,n-L�B�S(�]��%�]�NL���w�݁��O:!)Q1�;��(�w�yQ���Ė��Z�����A�"!J2֕;������:t�����)ɯ�e�Ŏk�e������y���������/��g�GC���?L�~��� T8e���7H��	�����Do�QK�������UA� bq��J�Z��'�O�� � 0�� �)��p�j�J�6���X���qV8*-�uK0��XF81��TamXq��������}�F��A�	"By���ڎ<���Q�H.�_$�4�P�� �Yz<�����J��S}�����h��<���4�i�X'Ÿ&ĉ��w��D��;�7����,k �֢�EN;LzҢ̧��v6S�B'�l���Rwӓ}C��pЏ��0�כ' ��j*T/�z�b�� �K���EJI&*1Ɯ W�H�dVHR��l� ��K�^��S*#�}�:��'�u����H�n��clí]kϩ<���&Y9�C)""�r �o"�a�jt7I!,�0Gץ6��A}r��^\�PTW�Ȓ�qI@r)�ApcjIb�!l}3� �yf
��E����lڑ�� �e�����@FÛ��_� �XS܋��A@�i+����K�1�SV8w��ݢ���Ev-1��]B�\"� ��%1�q�@��B����d�E��1�!�w���U��N��gҬeK� ��EsZ<�tN(ה��W�U Y6�Fth�>놎8�M��f�j��Ye0E-M0�Z�;��,�[" ;��Oܙx��A�UdH\�����0�QR� 2v^VF D��3� #cy7MQ�s7�Ca��@D�B��XM	�8��Id8cϨe��^��PiYeW� ��Z���b��س���d|�2#�7�L�X0��:��Cէɚ:9U��p�$�L_+8�d��"���\q�์Pֹ�! s�;a�u{�@���N�6�d6eAcm�nd�7�#��xc@|�yz��,P� 0��@���6�r��amdl0a��\�X�H,zȴG4��41"��۹��'�G*�81?Seӑ_Q��c&='�a�Z &��Ne4�ΰr)��IY��t��MB�\����Hܶ�|�`�I]Ks�el��@�'��y�E�c[�ۑ�E��@&<$dg��.;��g$4�^L����hK�i�>%�[�]I%`�-ޣ�8�{�9�G,�!�A�����R�<sR=3�}u\U�D��0�Hn�T
��d�t�1�'�cF ꦞ����8p*�RwI0B�\Q��&X-�X�`u��d)┽D�ɘ�Yм��;3�&���?H����s�dT����R�hG��pE�Yi���a%_v��d-~l�ך�cQe�$[F�##"Z [��V�m\����wXE��^\��O���/�����M��싻��d���� E_�+��$�B��A
�DR����z��wӽȁP�2���	�J�p�s\�]�2��;�����I�n[�4�7-���E,=ܪƶfI �B^n��������<���󙑎�`��un������V��Ѷ�_|v
�R|]$I{�4���L���/u�Z)*1Acb�[���2b��k�ʷů������|���qH��q	4j1D�<�Š	} ]jB�6�s	T5�K��kW�Q`��wn��o�Ȩ���DbEI�������k\���P[\��v�G�\�Q�+��u�Q�,Tcd���-[m����i$I�* Ť�i��ck�K\��k��;W���\��b�J�6�o�ќ�kx�k�_������ƮZ*�-A���ݮXѼ���K�}�T����t��ʶ
��*+˃��ܯ5rۻ�+y�o+W��LI��m���5%��;Z�r�v�r�W]��5���Z�E}��W�nZ�U�]��X�폶�B�L� �DD$�QX*ú�X��j�Uo�k��儱�T����M��6**)�Mb"ض
LX�bű�RmF���"�I���]�O��g���1A�5g��uh��gus����lksj�EEW6�k��BW��r��O�w������Ԟ��������l����e�����[�����A��[�������PLu�cm���K�\u����@��ՙ��M��k��2j���d7�$$$S�����6�r�ۿ;��'˻\6Ѥ���.#/�KEjT[FBBE��t�4V�\���������Dcv��Q�p��4h,A%D��ȉ����eʗ�I�A�0�T�B�C�A2Dj5�m�͒ƊM^W4�ƍi�nmQiwsk����)�˖$�ڹ�}�+k����W	tF���R��S	Cb��Ey�EXű��*�J�H# 6�2�A[��I���7+t�a4DW���ͷwN��˛Q�s���k���\�yZ��1�G���v6��V+&�(����չQh�6�.kV����(,lUh�*���4[Q\��VܭW�u�E�湢�w_撌E�웛�I��ěTm��y�^m����\ھ{�j��\��βP`J1W���j,@`�(��k_�5\*�-����2����wv�Bs�0_�J(ԔA��>+��wn{��W/��-�,Qh�ƭ�^\RR(/+r�1���Ouͼ��z�,Tj5^Vū[��	;�]�(���ut��0iݼ��b�W�sh�D[�܍�Z5�t�[�k�j��W�5�D\�\�s���C(�.�����s&"�k⫔W�W5��V*��^j,mo��ʮm��kf��[�n��75s�5^��'8�f�Cd�&Ɗ�-[纬j�RBDj!tKD@.�2(H�#���ͫ�yn\��wv�wu�\��"�fP�tE|U�D�m_��.���T�*]B�.��T���׻��n^k���\�(2|릞�k.j�j5ͭ�U͵�mn�4o7QQ'ǖM头����S�q1�p�Q�v�np��%�	�B	.�6�tF�R�����{�����ܣE��"�-��!��;ww3���d^]/;"F��Y��*�j�nm\�V�Q���^[y�%�n��mt-A�$^ouגtl-���1�"��\�v����c�n�k��"LX�.O.]�K��Db61o-�A����TJ��ڴڮ�|U�9Q\,X��ڼ��K2g
�T\�8Q�{�R=�[�����q�#Wuؾ5\ؼ�[�-�Z��+W��_V�������lh���W��s^\�=ur��<��ݹ���4�'v�&��Ca+��[��Lh�r��[^iJ��Z�	h��P��	���^V᫖�k��Us�v1nQr�뻮���7)�1<��n\���,y��#��	�\X0"�"H#t@��-�-k6����o+�cr�h��I_J�$�n��X�Q�IF"�{�e>.����˸�<L�w/���wFёΎ\Jgs��4m���mV�[�y��ncZ�k����m^wN�幷J���n�L�Mҹ���f�A�>w�˯��H��{�ț�]�d�8�V+o��֮z ���Z
+�@RȖ��B�ސWwN�ŴU���t[;��`�|��M󫕾5�)(�i\��a(������z��t��vWk�HN����h��br�1sr�wk�F��m�Z�m[+Km�⳺���msnr��+���|y���wu{���[��!�`Nr�sk�堌{���#�Nn��/^q=�L|�;tJ>N���5��|p��|�O��F��z�P��� H�x_$F�5����w7+��b�S���\9\�I�u�.]QL˛��	�bJl�n�ƺ
J4��,��vs�P"�ܩ�����$�� � ���EBFD��e�}�iS3K,EDd���$f($VDr�@9��ң���w���<b|"&�p�H�_h@u�v޷�5�vu�uj��x��� x._���쿟��#�?c�_��$�P��7�%�����}U?�'�[�����4������6��kO�(?������?d*y�vU�d��ҋ�G'� ����4IE���|�X^�$^� ���`�����4\u���B��Q�r�ڀ=+M�3�bv���hF�"�4�>�?��R�{��EE������/��q��+T��/�����V~��h��=��9Dɘ����[r���:n���
�vk��<=|��`%�ӂ�x?���v&%�)IM��=�Ӵ[-��D�1��g��*�ؼ���;|�y���%`	�z���뿔�6�̶�	�/�Y��g��/:��M�D2�!&<�\/�'�ī����3��-T�Ԍ�W2Η�J�m�I�?���t�4
g8���V�!���zu݂�Qhr��2u��^K�Nq�q!JD�Z6O�Y�闋ة�$��'��Ӵ	�}���I.�>8����i����n�Ħic1�6-;\ר�^NwF���Z���r��v���4��{|puw����%�^	��N��EN�86җ��
<Hp �[�a����Nb�����W����z�ΐ(�|^m;��gB�vA�y	+�W�I?;v�	�g�8�'+=Fs��(��[�T��6�Bo7s���1<rۙ��Q����ΨT�dw���&{-�YTA�Nr�q�z'ů�� �r⿈�Η��������4�]A��QY�z�|Ys0�
/��=�����(9���Ѡj���WCI:R�W>Yn�r�Y6�/g��,n�;��Qk�1,Ư�N�M�`N×����o�2"U�C�Z�'���P��^Vҭ�.�d�
��5o���*�%.���)��r�,��l|�ª�ZW�!����j��� ��3�SK�j�ɏ�p�z�"cq)s�B�:ɅŶ��6L��Se��C�"�N�^ԫ�T�d�gl��*��]CU�d'Nw\���OM1<�_Nr�C4Ю���\jѪ�k���-2q��U�N���&�GR��=j�4�¤,5��~�β�*�<��h��9�pC��r�>:����Hٺ�����0�W#��1d57����Ƀ��K�94���F�8���>�V�V^�O��3��۔��.V,��MĈ�d��wZ^~��/��݈�r�6u�W�E�B�-�_R����d�V�/��O�����?gIj�%����]k=�L��asf�[�*�{��C�b�J��Q�1+<�e�����瘑��W�$l�b����{6��)h�����ǔ�^��FV7{�4�b`A�V��Xv*�u�J�}j�iQ�s!�¦��2`�y�Ϛ
v�t�
^�[!�W�M�#�r��[�`��č����5i��ſc�5!&@,F�K��[H���zw�FR=�і[A��8��^�l�x��|�����[�H��M��P&�N�i���d��L=Šn�8K���]�Se���?��L;m�=�(�u���Ht�՛�t�s�*��~H(�:�4B���~.�ۭ1�������T�F��ٗQ�	�����V7�?#�G��fd]?����=t�M.ٕ�Vw�z\���U�HNv^�)+��WE�.ѕz"?�	��Lʦ;��曚ۍw.��ǢV�)�w�䩣��~�&"1ǄM���ԉ��Q�0���}�;U'�tU�(��:�L���>W��<@ �9�{�9�����齺,�6�}mv�d$`� �M�e�h�2�f��g����E�Bs�;쪛л�s��ub�J�y<�!@w-M�!cê(��\N�����	�c��a�l�~��"������A�l&��G�#<��Z��c6�/q*PY>q+�.�E$���efac�����J� �.w�#)�^�x3����^Z��`Kᖢfm�d�����	t�Km`b7�2��0��'aeԔ秊;�Dy���V��)����O��P��(0��+��%��6]%X
����wj�7Z0�h�l8�!��xN�t��H3T�a�M��O�ҿ� ?]�u���a�r��K��X���O+��_�B�Óφ}���>q�RF~�G�"&7���Jv8<t���X��$'���XQ�XM�3���S%�Ky`=��9�![wO`���~�h~�@�����~Ȫ4�+�KM(7������҂RO<#̪��@I��`X'�_���M� t00��}��U�����ġ�q��hO�"�ϳB�l���/��$7*Ҁ	ɸk�}A[��~��eӘaȊ��R#��)���sJ@h0��~�(�M4s��%>�1"���I���ѷ�E�	{��:��1$�lo�Z7,� =�lT;6k����N2��k���eq��=�9SrK� �j*@aw�ǂġ�!�]=`z)�yZl���
�����䪷��9�%7�+W�	I�����V�B��8��<5��0�����{��P�\�ۈTd�c��KДB,�R���!r+�6/F�>|[&���Jz�j���1Ey�8_����z����a�l��縈*[�[�L�P@
8,$�G���(����D�4Q�K(���!*p��`�-D�H��0�A��5I����__�C�i�ukma��$8���'�c68��l���ܓ�$�Z� !qH�Wv��!abr=4�/6ab%&6���θà L� �﩮�B�98�8VN6b��*�F]IA/���Pr�)z��@�dJ��m��S�H��ɥX�-�Lq�n��mBm2&
��V��iAH�m���!
N5�o�[0�,Y�Y��V�fNp-��D�|��	ýIF��.V�A�O�$��֞A���j�0I K@`�aMX]+��2��8�Q�r�I3�J�RأF��	!RS�)"*�eV����]vET��̒Dl�"R��q�q�^����w;a�vZ(�R��v^A�OAC��u���KfXه�?���q���;�;��'U�hȐ�Vd�Ɣ��̂EzN�yW��^���0��2IfČ`���kj ��WM̃4�p�iC�3��@��>RD�$�%�$��F��ńv4��#��e:=�]���d�KH��ft�'��Fզv������1�؟̩�J�r�f��McN��nQ�� �E}�����?e�1���e��Y}`޿�Z� � J w���VA�K�����_���?T���>W�I]��-3%�X,��%jKg�*V��M%���I�R�ji��h�(ƒ�li2eU�'����}O��~N�G�~}PW������]���p��� �kclU�[U��V��P
��� ("��B�y�^���<U��W]�t~����ǫ<oAߺ��k�<����d������˲W�8~Њ��������O�?-�?$��o�'��,1~o�$&��/޴�Y$���2��q@��+�R>s����4f�n%����x���1�e&�3�Iq��%b�E� �[�z���7��ks�{ABƇ~�H�>��7����]9g/�-��{`��v�M���#=�5S�'V��:�M��T:鬏u��O�Y������td����7i~��Ǯ�m�ea��S�̼�	�������c��8��2�[�"!�]x[A��V�H���ȅې���Η��#�.s���\ﻝD"@��N�!f�cO3ʤ��#���=\�5Br���E��Kݲ�1\F�jub��w��Gb�W�~�r�_@w�M�,��	�Mˊe���A_�zi]�}mwIqz�#�O%��E�:�ɣPW7{lӹ�*|�/.�'CO�WRD��(5ގO(��o"�$�1�U��#�t�\z�W��D~�S��4
{���~��ƃ��uf��$�&��9��[��7(��4���_	o\ }������'��z�-M�z����A��Eϼ�����. azɒ:ov��}<'��Sy����2^�t^o����Yu�9ps~H�*��A;\��)h`[r�`�BI���TH3�IiQ-�%��f�W �x6�+�̵�Y�x4�|�!�m��S|����&��<�Py{|R'8z�j��}�j�*�+U��9=np�)뤩
 �A잒����h���b�`9h�Y"uO�[���J#�aPQ}"�6	(�fG%�JD�rzz)���E��*J��冻s��FO0d�3y���ƶ�<��^J�a)�D��D+���:�oÇ�u��d;ɐ�S����;x����#�:���	�uw��kǙI�y	j���C;Gtq�i�I;�Vya����Z��&���O֔Ä�����0�7�2w8���ۡ��Ʃ�^6B9�E���pm�v�����ys��{Q􏍵�Xf�]�E�)}��!���sÆ�,ՏC �n�s��α�����X�{c7�`3G�(�v"i9�D�$�^��`
�T���7�5�X����Z8Pl�L�~O�pU��Gih=RQ���^Ajc�~z���2�n|;���y!���c��ΐG�?¡�ל�zH��F�I�+}V;�u�؝��,� �̓{�DH�Z�9l�>��k�n�[�Kf*X.Y���mCI��>�1V޵���BeN~�;z�g�Km�z��l�y8@k�7���4��s�U%�A�j�cJ��Y��+��8d�Pɸ�jw� n.P*���ۺ51_�H���51"�Nj����)-|��S�}�Q%w.��6~QV&~������7��6����"�&ȄM��iͧr����JtW���	^���%{'ӦP��4I	�ß�t���m��G�ꌂY��!'�X���>^*^]���3��|�pm��W�ʣ �,�'�%�v�r��<h/%��cDs����r�K(U�d�\3�t[�Dy��0��
M��Q�xy�<�����p�x�+�NW�F�@��4��l���ct�x�7�j�+��T�9ң���i�_=�H-�
/H���Zu�S�n���<&VԂ�p�dpF{�+���F�6��?nNUu�|A�툯�з�~n��Wї-j�A$�|:Rp���vn�a?QNdU8:^����;_�0J�%
X�=2��T<FJ�H
�i�B�u��l�O���R+�=���
'��)}G��"[�Y�շ�u{P$=tP��s����a=1\��G��=E�S���K�Ky�+q���>��}2B.��Q��LioB�RV��b��j<wP_҄s�!�v*
����d���LX}�s�K�&
5�x�_�����ko(�W�сo��d�r�.9(͌�5��kA��'n����vV�~^���'*-xɾݧ71��ȀwuuT���S�o��]E�N�H!���YI�ü��a&4O�9�9=�؆nc��q�o%i�����ݾϗ=�����g�V����_�cm7�?����?����tҶ'q<�����'Vkˁѹ����;��g���}]��G�����������g���?�����E��)q�4�<��K�����?��w�}�������(���i��R��ӌ�@�r?�`�(���I
 ���G$�ɐt�ʋ�<�_�I���9��8$�:�@����*���,������i��Qy�"����v����j�#i�ޑ�Wx*4�L���gJ�y�2R�p� ���Y#QQC���R�����HB�N:�لf�]Y�}2�8�$��T���q�u�����0�\t�!�c�-�Е�P\�� �j�Y�
M��)��addIe A6����4g�xS�Y�`X ��U�A+����y�"ĕ��a=��Zp�C1�r��+�D���$�e ���CL����Z�h*��0�JYֿ*�8.@Brc*f����OaF6�0��L����0�M0��KHZ#�!(��x�3@ڑI�j�&d�	��Ka��U34�&�b�M@ޕ�Ѕ�Ra���Ie	�-B�*z�&�]W�
���-�o����Aׯ(��\���$B�G?4� �ʪ2	9�:B���N�M��h/<7�c%�3趼(�k����H�%�V�ߒK4QO݆��6>�Ev.)��Od+�E�@��A����X�)�Z�ʘ� eN��8$�{$���<L�!d0HYh���<��a�V�b�0���l�pu~�̸ˏY� Tc�1�t��Ip�!��kp��m��j��R�����F�G$��eٔ��NJ����.�y��ծ�L20.@�r����2 ����N�Faa���S�W�a�Kh��O��q��N&3j��,�p��<qEFN�^��H��%�Xcm7Hs����#EؐEP=$������-9�rR\*@Û��W��Z�I��'
�#��rV�G�<�m�bN���t3`�s
X�� ����P��q�����6 pDPJW�	Ǣ�F�[����Ĵ�� �jd��&Kh" iB@## � &�C�>�[���>���"j WpPCXP$FTD�$."�*4�- �`,F�Q��`{}d~G������8g���{��������+��	�@/�~/��}�����+�}�1�Q�F���b�8��i��Y8�����|������5;Mye�*�����_%����`R��^�J������`  {	`���so'�>�x<vI�?�fY����Н�cVX�8���ڙ3TR2~�t{Ly"i��*���!�)W:|e�����I-�e���#o(��!Ky,[:U���*��?�T��%�g!��E�`�=��   B  � �` ͫ|����s��7�c���=���(�*�,���-/s� X���:ۿ�jo� q�=ۖ��*mj>��zTH������-����ׯ[��:� �9	�v��1�{)îo��֗�O�+~=%�1O��cA�@����M�D$I�l>�;9�+5RΦc-�Z�֥���-M���FTK�Y ��4:�Ć������+V���&�lƎ�o��������Ơ��g��{{�yS�� w>�����o�}�/��ź��Y�j*���Y�׈�����wS�;�a��C�Q�4�H�G�W,d�r�	5�7,�.��ic$��o�rj*�K|v�z�&,X��xd�k�2��te|�Ow������ͱ����g^�#����]��+h�&"x��o���?&.�w��<�lա�;1h�N�k���|Ԑ�� �A�&��Fqi=	��,�O��T-zf�[��G�).$����S�2����s�ԍ*��K�%��Vr�gb�=[M��F��&�Zy &~���C*cU�ˆf������(I�Q�6��1ԍF���2�Ǡ�s�����y٬WR�E�"��:��^�#!)�Sw�W�P;D֩.F��f�@ʤx-«JoA�D����KJ��<)Sv�of�;ivPqdW�p�n�M��� QW,���_N�u>��˿�K�q�#��'P*u���<<�߬|�A"�P������:��U�Q�ͨ��G��(Rh�2,��QS@����ڶvYu'[�R�xC���5�c�䔼��"�n�'̚V�[ѭ|o����K�������5�gb+�i���)���+�0� z�G6N�>��L~^D�-y�y���7�c�B�^�=��ruJ�;E�-�T�<-J#�f҂/0\"`��և�����9��ǕʺCUnh���-�)��.�Q��\Z\]��+��Vt�� *��م���2��qC-7}&D�cMv��{�����\Z!z�/4�=A�oD��az3��R��ʸ)�P���c��<ݿ�ۭ�3X����ƞ1\�N�q��$��z��CE�d&�W/�Rv�����/<}�ڛd���a�3�v����f��@s[��<n��%��i�^���ֈ/eZ	��l7D+�-��n�ȝ^7~�~z�̔����#v������^oSc�{z�yD�I`�R�o6p��ς^;;���!�^�s�rx.�q�����RtB�Pj�l�p��L
'�/��'�AUJ\om���0��Q̓΃�ʓ�_�#�3� Յ�]8婻%sN'�(���Kܹ?�]q�t@P���hKC�{�3Ȣ�&5���<��G�T�r�l|��E,c��z�K���X�X����T�S4.�c0�&/Y���g��l�Q��{�{de���m�Ί/�JP���W����7b|�v�ħA����C�wxm��"�{'״�n.�]�6yJv4�S[��f�-^��Jj�!�-z�6P��Cib`(��ڌ�ƻ_�s�(�����B����U���ޢw���P"L����R�'BxP2f�������*��i\o�&�ct:rp�"�d�`��v>�.��D���Qa�r((q$A����︮M��z�9}���v�>���:<X��}A�uR�c��W,w"=��ܽo�d��^T@8�(�F��[�aKཞ��޹����b�_<M�M#�L8�2�C)����U֋��(��b�'�o��0>�	Wä�/�H���x��$�{��Q��0����#;I=��Lw�?��3%n���M~;u���w79^kv��H�Eb!H� `�U��x΃���>��u]'M�m�]��r�� ��|���9�}�z�<R��$A�a��K\��Lt�@%�U�ahŊ=p���� ��Se2	hRNK�}O����/
�R�A�@B��Y��Yu`9#�!1(%e�|�Qq@Q] �v���5	��%�V�_���Т��T`
hu�h�WI��^�O��O��q���ZV<�_ܬ���R��]�ht�}��{2�J4�UPA�$�i��i�DH��vL��QP�Mxa_���ɝP��M�'*��8c���f����LK�-3�Q4����� ��~�+BYY7'ZǊm�,���I励s�)���h��9��V;r��.��:�Ch`�"N;e^U�x���j��!���H��jtM. �Z�m��&+*0�%E�����Z�xɰ�YI�d֠�" �U'�7�rށ2`Y�Oasep�#=�`�W��XTK{��N#Q-<�ȭ��I�J:��nq�q�!"Ma4�8Ƌ� ��!��9��p�l�MܝW-����<x���|�ik�6�����GŻ�))8�O:�P5�6%�HI[��UҚ$%l��n,mH8��$2f�Q$�}7M �"*	�QF�� ��\I��Tr)q�F�`,�D�I$� #$���΁�d�ǅ��1x�ma�9L�WR��N�d>�>H�՟�0E�(bBp�1���)c��L��N	��/0�)ց��d�{U�$ZPi,TM�Y�+̸�JV��pB�n�Zd�
����"�$��b����G���fz�.������E�­x�JV��DR.nP0�N<dIQ�> �M�N��%�x�I�a��/��JJ'(5kWe�0�l��Pe��QF	�A&BA�9\���u�mg<K0��`���,@�)�p��(��6�+��jd��a6���죤+�Ŋ�p�D��H��\b�5,jeHֈ�5���h茶�������[�!H xN���������<7K�s|U��_���{�Ro�����.��������F�S�3���"��P"���i>��K���O�E_�]�$��1����&�(��R�4Г`��b�>ȳm��mS�5}�/�\��H>�$/2�R�k+�y�G}5i���(2�^ӹ<(��q�����H��0utlo�(�x�+�>I�q�$���1��\����2���|��7.p;��Y�4ई�MQ��i�����c��G*��q�#��ܿOw�`��P�(�W�-]�>�k%���@^@�N�P��=[<{�ޓ�g��{9���w{+��ԻJ!?]�n�d�����^T(L�J
�G�ȮǠ�����S���/����rl��Vvhމ��լK6��I�z�"�E�Q����Uy���K[�r��|�"̦O���X_��J3W��ʇ*�/�r*�^!}0�$X�:6��馰���ǅ�a�9�G%�N��R�j|�3�e�t�(��H{���ʘ�m�����*���d���SH���7��w��9-;^�;�Vo�o�I�Z4���2m��l���D.��uK����8��'��7�F�w��/&g���چ+t��;�yC���
����{f<��m�+WN��Z`�}+~־Gk�?��[ɼ�M��%�+/s�-��s�֭ܵ5p�7	�TH��)u��w��=2t��_�S)����4r�Y�[H�]喭f6�yq�%�y��4�5R$<A�q�W!����a�?B��1�����:=�I|Ǥ\��'VJG��nr�;�:�<8����5�o�|��i�Iݏ�p���n��0���;��6Mw��$;��rz�=J��V��W�������ZȞ[A0����l���S~�*�׏T��!W��͏��V�������*&s8��%�g ��t˄a)"��r��r3`C���[䍝<T|{��_&�Pb��>�V�U��O$f&���ư��uQ7�U�w�s�7�J�d%5�%�5�e�tߧA��s���Ke=��bxʨK���AWxjl��1J0h��Y���y%�D�[�S�,�R`�=�5�C��5�0Ǽ�M�%_���}�T��eF�&�]!��%��d�F=�R^�Dv��?��dsξ��zsřt�^.6�e��G�%X��K��˖��㦫U���� ��9y<��3w%�T.~c
��Oȓ�������뇇j;����zVM���$t��Z4a�]��	\���;f�]��X�$B��g�#9�AY3�X���2HŅ��/ܷ�PEg:fEy}à�����y����u׶(~t�2rQV�:�w4tMv6�p[�P2M��:�����ܷmmꐜ�L�krɞ|Ns�+��3���N�zÒ�����V����b� �~�bd�7���/�=}o���E%�=�A+P��$f3w?QL؆"�E�f'E,G�;B����Th��ʑ;���B"u��&�
/1��V�>xN�B�^g���!޵w�/��L�`�>�y�^T�k�k���9#������&B�Z-)��# �w2J$~���=��=b�|�����9n�sAz��/T=D����%��o��`v��eI)�J
�3��T����Q��Rso#��N�[ǌ~N��W~<�Ӓ�l�s\̢aI<�Q�V��2GOL�+��~�ҽً�Q�7��r����9=%&���s+�-j�Lp�#�������U�h�X!��"�$~�����i#J|�Ƈ�Sq��X��KO	���Yl=U�iT���a��'u��x*��N˫��bf[�϶�ST�=��\���%������"``h��kx��q��3a�}\%�RJ\�9���d�h�Y���עJ�1|(������(�@U�/��塊-]�FBQƽJ�=�'ի���y��.��L�����7�m9��
�5+x�z�O�+*|�K�y��z�+J�Pb�����<�J8������<~�>=u�	�+mE8�.UAY#�R�.�Op�����d�#�������x>�?�7�|���D�������dV���eK���c�@�O����E��Qi����-/���?��S�{���._8�2c���<3_��j��u�����9���������[���k�3�&��H�u'�2�b#�	N�l$��Ҫ�L��huM�w�M�*�B�t5PT{SFb�RdȂg0Ⱦħ��*|��Lx���X�iG�f����>������U����﷎�������eXڙ  �AXʥ:+$���h��m�z�@S�I� �"9�Д���¸�p"�J��T�'�A��K�% LR*2�4	�	T0���U���}�hJ��x�D�Y�Nl�� �R-�$H`� AS��z$��F(n2,J<&2qjq��e�0�ձ6(0��YW�P�����ap�r�*p�|`�&F��&Y��1N�p�=-B�H5O����
E|p�A��?���0��z��2_� ,3~Z9#�lm�>�Li�!F�S,��9B
<�KRQy�P$t�"��4b�d%�9����"@\&%�}��i�j�Џe `�Yi�&!z���TM��ng+���B��h��EJ���-G�Hf�HO�U��)o��9����[F>aLj������Ey��4�`��<3�K�Z��횘�����d���������4�V�L��/�ҝ�ʂ0 T	��))d��ըu

P�4g��G-�`jg�9�(��9*>��&&[R1'-��D�#ҋt����O
���ԒR0ʌi� ��'����� <ا E9Z�g�DV]��"�g
AY
H�е��2,�����/S��o .]֮�`#�* ة (w��:��hƦd��
�j�X��4 �I�$� �BF��_����+�_G�������Q����������/�����)���$D�!J)�?�U�&�V�W���`sݹ�qKMy��%�S�f�<An�����Um9����42�4h������������7�/�@���qW�3���"^t��Û����5x��(���Zffo^�Z ��O ���s{F�©i�f�$v�I��Nk�[԰	޿S�\]���TC�(��6j��b��[u(����ފ�S�Fw�B�{�	�H��/n��F�i�.����k=y�3˄]{ Mo���ó��&�Q�hᚭ4����*-\�к4t��l����J4���ފ�����SsA�9E��Y�/�)�̥]�%��M�6)t����Ū��;wY��3�HB34������6�Z����"V�6�εr0L�U�f+�&+r�ߝ�Z�2�����s��fs�hUW�n;��8�F�Ψ�ɼ��P�i7�ގ��q�F`��"g)f����R�c��#{����˻�p�^�_ %q�N{n���<OQ��{$��zx��RÓX�cB� ��C�G�o1؞��"L�{�X���ֶ+�v�]\�0D���^���D(ʳ��_(��L}�*#�{ ���{__�I�B������?[���}�_T�~F_h��~B"A�y}��qY/��%����D�H���e�����d���Z��ߨؾ�M���߈�Ƌ���_�
Q��`�럗�S'�9{  �2��)�o��+����'/s�!�BlT,��Y&	r��7Gf�Ko�7�s�A��kE�Vr��Q�nc;� ?�����i�^���y�ʇ��I���t�;�I���*
E=�
���[gcM�|�P�g����`�!;��&���O�Q�9�8qҸ$V�V��_�Үx���>������3�B��j5;z7�P�T+F)��K����&�p<�b�]w��_˧`�#�r�u/�o�P�6F��!Lc�� h���c�щ!SF�`T�vt����U�i>�'T2y�����1��DZE���X�Q�N���ԉ�2�����mY�y�g.����� �{�d#�k��B���	�0�9�8�\b.rTO�ǹ;"ڙ�ɐ(�JHu�I���k�lSo�Zf��.(UBs/f�!�:t˿=��tqz��l���n�O����ȺL��,�$Gn��0y'�;*"+�z�H�㎍X���"�;ʷ�q33���|L�c)F'�[-�ߞX�)k3Lp�t*��޶S�q�D񩮟3� �UӋ2�>1�������%7/��J��4���hXؙ#(6֢,��ϯ�%����Ӫ�à�mb�O�.T���-U@�h��TM�u�a�匷���S�Wxu�Ή������з~s�׌c���I���x�1��^~Ax>���+P���]���QW��k<���~^+��i�j�@�Y����o$��� ��
�T �^���(�)�XB�LLJ�tжH<vk~	�7��v�ߵ];���t�	
�k�!]T�|
�<�A�y13'��4��µ$PM�yU��WB�\�A�ǚʯ!���:�V�t,NUV����#zJ�sc�Ǹ�I����P� ����Dɱ�u`�4,�#��U���1�< y����N�QƮ���_nVk/��z�E��b��Eƶ<�Ȼ*�%sV�l�z���/������p08��5�	�d|�����p�	�e�fL�of���^�q|��BXg���6:]�+���<�2=�����b�C�����i�|�͂D�{Sf��Ŏ$)Or[G$u����O[y��Ҋ��>+Z��?C&�t9�X|�r=��+�1�x}���j���!�w����W�A�̜I~����3Ѽ���ϡݒ3;��I���i�q�M=�1�_�cHv�Fv|drj����wy��zu��g�%e��-C<�bz[��:�)�����;��(��wc�9_�z�Gq��pr�������e���$��y���栌<=i�)�5lp�[�^�O�nd�U�2�u�U�����}���v�E�Y�=Z�I� �8�8�s	��OASx�V��}�^a��/x3�C�F$�X���,٪�5v��,3�ۄ�*|���)U���L���ԙ_��s�S�M��P�H0c�6~zD-��u:���6�HL.x�2(�Z�z{kA��xv�ϧ�Ζ�	�/��?}�:5�et4=P�^�,��Fg��/���% '��� 2k�I��/�`�cK�e���i�°�Ce�U�Y^Y	��c�^��у����_-RMǢRE��\b!�^��%�:^j̻�e����S#�y��>&�t�4�#;0(���,S��Dϸ=r=q&C��!�V&�n�{e�E1�^;B��뙅[,�9̜S��K�*��P���bL1LHQ�zw��M�ȡ��ט�i�Y��_-�GS��w,�k�4\��$�>��:$<���_9⑙(o&5�Xw��<��*�<f�f9�W{���Y�;P�Mқe�R	�+�E�-�D��6�\��w�h��<,�/��(Y��VW��l-�G�HQ�k�����+м���j����2���u�{����?�����F�诵���a���Dϥ�>���T>7�Ld�/��KC�}A�,P{�4)
2'�#ǿ�z��2�O���|J����_���M����5�M��f���m�q�f�����'�ֿ��.1��4���k<�p�ڌ��^�5�pIT���-�M5� ��I�52����H�dg$��h
�-�)����D*��X(��`a<��\rTP��,a�4F�Zhޝ6�D�M1�-�5�B��+�.A
�@(� Ѓ�b�*Bh�H�P��J|�$iӅu�]��
��+�΄��|�f/���?�������?$W�ؾe��|��T�p�������ʒ�INy2?+�.�
 ���q���$��Ȱf=qe^	�\y�p	2�83��(��(E�&0�W��|x%dE%�!��qQ��V"(RA�8	,#�
;�o�V�CoWkC���c�6�o)�-���/��X[��g]O��V������������b���9�Ƙ}�I�1QP��bI!$�ʚ�� �x�����!:>� �)���H��,�>�e(�Qrl��@��5@'��ߴ>>�4�ZQ�Ei��Mch�^��q�m���(��$ �l��1�IU8�(�P��f�D��DVr��ArI�S٘Ǉ-Y���䌳1��8T� [*rG�)���2ƊyS��gF8��$����FX�$q��d1x��ҏ�<�>���{v��eۿ������|�o�"�P������$�����DH�0	BIAah�l�PSS���ʪ��=�x�w��x�2"=�T����~�־���_m�5&5�V�`F7��og�s"��ܺ�S����қ��Ѓ������ډ˗��h���"oDMWB�틺��C��80����W����8�-҉��c^IXC�];39�ڤص��<���A�Ǫ�z7������=���_:��50��2r�Α�e�}��%c8�Qw�U��A�����c�@��`[X�vΛ�vWJ��Ҩs�ٷ�S���sھ{�G\\�����i� �w4DNb�u���v)�mJ�wӂ��b���|w �	-TE۵��͊9�a�n����O�WH���ڞB�"��aGt�!&]ӫ3�ʂ%�K�wL�h0��(;55DY,��c*iR��q�Z�j�:aF˻�#��5��a7၇{Ne�quW|�$��Q/	��ZPָ;�3af^vZ�}�}�Ͼץ����ǹE&�(�ӛ@���'�p�M�g��Œ��+��g������Ѻ.�V�8P�6�hҳx���Wy̈�S��K٭\lq���V��w�TڬP_�6�r�{�!�w3�\T�*��ɵ
z�&(U���rAudf��sQ)Y!�q��+͗�X�3�5�՚���1Vf�Uw��ؑ����l� +aQz@�K��x�uf�JM�;q1�Y:�9��3Υ�3�2D�.�S<��X��S��cbtR{y�E�8�.zJeĒ|�v�p���|�J�.8�P�z֝��,�%���	ӱ;5�[��v�P"bt�˹'�DӖ2y�����v�V�����(sx?1�(�(]�f3G�k�ݩ�(�&�+ةD-������`�3�0;u���G��4zpBT��\�
�$�$�Q����?{���1�?����k��6w�S���8�G�|�����|�~ID�?�(>8���#�D?�A�߅���BU�4���?�|3��0��~�2G��EX��{"&��v��vW=����(Q�`{{l�_<L~��KeZI�
y�V�V+���_I;VL�:��&��!�p#~gG�q��9���ⷚq�?�e3��1ΐ-��������D�g�GID��7y�ȣT�{t�d���[�:�9qn0�����Q$��n.ً�6�}_ PԹ  �����S��?�j��pÜp�&��̆�;M�2x�x]������N��J�#��<K�3{!B3�I�;#X�\��bb��#���lW�.cr6v�R��U9@e�sf��'yո�b��u��t]8η0�vlz��˩2Ȳ����UY@���R��iwos4f�q�	�kOPq��3ـ,	1d�@�Ua@�d4��vj3)��-T��GX�L��>w�O�tk��Ľ��Rc>�k��.��L*J6�_4wB���ݽ�*�F�ݮ��7b|wQV��������p�n����͂����v��-6�:?֖�� �%�iX<y���b���O�t�瘥^[^�s#�[��{[�8yᲱ�F���!�$��WĶ�y�6��nM�	��
�<����ɪ&��%�J�b�QiV�(����=�QN��x��ܢ�ƽ��nj��ĝ�O�?K�)����i%�{��cھkI�������[v�B�j�VN�>hU��(��A��ô�7eo��cF��{oD@�{uG�;\��9��Lϋfy������<#v���a�v�_]���py����N�nd�ڷ���V����d\��_k�����n�ȣS�r�:��{i���yuN�ͩnon�֍��L���6b��A���L�Q"��sQ���Jz��A*G孇�X��KQu�^w�I��g~o�I�	Ъ�%���<x>�#��h�(�h������ h�:+E�q��z͸ɝ(F�6`|�ˤB�������W�Z*�P��M3N�M.���J�t0>u<�A�KA5P6�B7������I@cV��0LQ��nXEg�J&������|E��X���c�2�Li�x��q2+l8��.���k^����Í����;-O��)x�	%(q���3(l�V��'yPadI��*޻vC\�Q۔D�d�}d�,}�n���� ��o+��3�m�O)��|�_8��ŗN�V5$kNJj�t���]������'m�W3W���:�j�1-y���C2����9sĤ$ݾ-��dh�&u=!]_��M����^Yƚ�|�O<����#k�׉X��(=�1*��;W�d�u�F�:~��ѧ��@o�^��M‒�fƤ ��1E��	i�^f��~bUh�MNugu!˶}�%���B��>��a{�|k�N�X��|D$Z�V	���^U� �7.��D$�5Iğx���z�
�"�/�A�R��x�Њ�J�]�C��՞�Q�~^�K�Sp��rq�	b���?.zYz�ڲm�`d�r�~�����|n-�0q^ć�P~�D�8��G>Ӕ�"�m�u!�v�"��m�I���«�
;�"'�����`��v��8�{�]�7?T���S�>�k{��mS��L�T��QK3D��ea4���PK����V��]Ϝ��&xq�{�s|�%؍A]n11�uh�!� ��u��q��^�������P�03��E��7G�i�Sr5uZ�ߙJT�����Թs��y�D��~M9|��]�o<�2���
��2
 �DHI���O�$��9��5md4�Z{��ۡ�Up�v���۲P��rf�S�Ю]��.aR#&��h��J�LwL}�(�;��2|����wG�{qZ�(O72��[#�ie{Ή�u|�9��j��N�Gp�y�Ⱥ�=O���ͮ�~�1� =�����K��(�	�O�8>_����Z"�_������XM�g���[����~����q%������۹����(��������������+[��Z��M#Ja����~��#���}~�����������w�G�����h��[E�Hh��1�rg�^-��X�tVR!tb@��9���e�3��!����x�9�oy�e��<q��7�q���#�&=��Ts���|��)�����Y��{��K�L��$���h�9֏d��%��9C�"�AK��^<}���'�o�ۏU?J�R���><|O�E禯ލ��AL�x	\ț�'G�	$6@�����L00IQ4�DĈ�*���B�j��ʌ��Yu#<h`|�օ`�)�!YĈ{-���{��{�q9<_�����گ\���O��v�1�����|5ޘ�[
�T�e]Cm��>}}���u�������z���˨+�>9��׌��1�4���v�й�������}=;�QX�C�}��������M��l��I�{W�����1���ˏK��޹]��3{�#y�k�{F|``ag�3� ���
|�h�G$m�#ˬ$E�@��8c ����>,�,��%��FBZ�@X��h�cd}�J4���cs�����V�֚�֓�����v�f`�=}�v�yo���m��TD�:�*J��c� ��``�����-uC�黦�����?O���ה�ZJ�����. K����/�ȆfQ22d��X"�T��"�Ab��_�s���=�Q9�E�v���|��ߺ��r����	>ʫ亳d|v�����|���h���Ґ��/��=?�?�r�����4���#nXa!x��(�����o`�� H���?C�f�D�����\.[��u�;w�W���\Dx�I-������F�Q�B���ƶJ ���N1��:�Y�k��\�myNc���d�є�_������+�m��}�]���p�m�ַ�@91�`<e�"�G�@¸�!�����}w�9z�q�s�0�
Qd�Fb�$_�?���9v��)]~�A2�6�:#�ǎ����k��!��C�$V�cr�T�t{�c�����+�Y��#�y���r���8C`��ozz{�Y%�8���X�S��:$�8#q46(��*V�Bm.��f�.4'�w�QϬh��ݏ����Х��E����ha�!:��Ұ*����l.�j�7��䑟�g��$l���}��L��wYg�n&��,"MX��\/!i?�lY���}5Ej��: 'P�z{��B���B��q����'��-�5�_�����doY�$�M]��fh~t̰!��d%�*��ޓ����v&�>�=G��)�bC07�E�C���q<	��eL&�^��=4R����#DքJBH�$�L;P�ƅ��tvѠ�ٱ���O�s&��+rVaw�|Ñ<��] g�N/Ω�tqyP�|%�Jz3"F0�~XV��F0uȎ��I��ܙ[�x�ѣ#���{��S�r�C�'xw�Ew�Gt�V����̸G��jM �0��0�d,
8���'U���Щژa52��{&�;�SH��?�V���7u��u��m�7�Sm��`Ԫ�[�Q*�M�d�Ƙ;>}"�����ێA���9��ۑWࡖ�F��"��pF���$K�A�zك:i�ڠ>8-�z�95w>I����5;#Ef?���<|+������U�+��ʽ��B����C��0���g�V��5x̜0�4]��D��aW��sx�}�X�d3�<����\�����-m ��_$g.R,fzJ��b[kk�ҹ�=�VeC��g��i�B󮀒���A���bo�#C�&y�G|EЃ{#چ.[�8P�t��d�̗�n�f��Zw1E��,�3��\���'�E�9���LX�H�O&4���1Om�9����[/x�v���i/����s��7�1���jF����KP˜����Q1Gc�Ɇ"J^�m��p��bX[�3��l�qH2�3TL.����;BM1�g���݋v�.p.��'�x�'<
�(�d����W�Wx���J�����G�^�F2	�.%�5z*u�{�g��NM�/U��G����p�,�IYL�9�r�����SE�d4��B��\�4��Z~��,���RG�VU؛Q��8Å����
hT�mm�Ju(�%��(�ll�(.� #�h�J�{w��S�-�n����d9�I���Ti *���}�mƠ�e9f|ܐ`���ԩ�w3K��:UvYJ��*<2Z�Ŏ*ɞ��F@��r^;7�U�}AU��'ҊlV&��=7Ԃ.���[���4�C7� !b �r޷��$���	���ŭ#���Q�qV::K�Eu8�{��:���U3�����Vc\����)�{�,"��#�9J�x�/bkd���A��J���,�i�SaP�k��l��w�a�K&��F��L��(�WU�zE�x��8��Y.�Q����Yv�:���!�KM��m:�&���]�7�$�ˀЇ{�;�⷗�N�;���T�Y�PJ]�������,VƢ��8��}��v�Bk/�]�U}i}�m^��F�M�\�mo�/��F!�g彽�l�>3l���ׇ�<\N빸�K�F������v={T]	�9����˸��Վ�q
Tb7���d)��v�䷺���t����O�˧�o��V����w]��P�Qb	`ABK:N^���m��=G�������O x��CO-�M����緲ێ������y�z��}����П����j�Q��{�ԟh���~Zp�|��4���_P�|������k�q������.|0��Ρ�>����α[o�hNW�N=O�}�w��;v���ސ���~�|V���lbw������7hmY��^8�;����u�W��_}�թ<<�,�������B7oq�U�l����{�a8�|K�}{y~�ꘖ�?�7LI����ĥx���N��p����W�?{[�կ��3�kF<�1���{{K��������P�N��3-
�슠�8z�2jŴkO�k��.2�.�x��0������W����.�-�2�Y|����|�p�ho��k�??ľ��;�������F�|��;�����.;g�?x�G��dח8�����'���״�3��sx���fzP�;74�u�mE�g���īA��v�w|��u�����^��ь8�����z5�sN����cߙ~/���ӵ<m���x���ϫ�;^�=uc���""� ���k��l���A� �� C�z/������]w��_`�54�2m�v���5�d��vS-���O���H��Xf�_mG+�����dT}���l{ӣҚ�F��_��)[q��w�f/�Ӆ=�p\����*g-#����U�two���A9�����u�]�|�b��d,��g̷;'���Ef�5�5T�Νs|VV��[�)��c�� ��/�E��ʍfu�ҍ�/��ca�q�ؕ�N�9�H�#taK	�ro�pڶ����w{u��;� �o�g.cNuGnm)�Y=g@Ν��; ��UGv����Sz���{"s.���E�G�U(pƵ�n����w]b9�ً�rl�(�pR� ��{���AQ���(�Jp��,\��Y70�:� �/�ML�����@F_T[�C����VY��"�x\^��{�yV^&oLq��)��eʄ�yv���R�]���5u�������8�;�3H������@Je���w;�p�F�93����n�y�ͩ�ج[��B5^�6/��YY;�2s�Z[B�H���os�*���L%"�b*�K����.�ov�<÷(�`;���nU��u�se����ս�2&�Q�ti=�Zɻ1uy�$�ŸZ]��ʑu��C�S��n����wK�EULmmN��C����Mj�ѷ]sr�ۼ:R�p&.�� �}\����5�� ԥ�����-ʼ���l=T�'����p�f�nUo{�g�v-j�rqڮ�<�*�4s3�wT�<�-1b�����	���=v�6�_�z����W*Lc�����%s��E�Ѕ�"*��mD�E��vD��O�v�z!gM8��j�屳md[�QΦ�L��/��)�ޔe�u!{7��c��trz��z\�Z:y5�U�ڝZ��gnr�R�5��s:ۊf��w7�uWh�`�f���5
��*E�:ۜ��7�s:%gn+�ˑFm�4B�j���<�ܛ��$���)S�y�	gK{�qJ��s��)���)I��1�x{I"�Vh����Y��ɶ�M�2�w��*kv�Z�'ncm\v�^(����嫡ɭ�6�,ݍ���.��w�iC�/��W�:��*��y�����S'��>�8=���)�"�fa�s;b�to[�u�EV���9��H�;pα���^��r�
%ݚ=wCm�Ruץb�ں:XC����0��Ʋ�j�����3��`�ʙCOS��o:5����{�B�{17�;mf��2�Ow
׹[�m�Ԏ�Q����}����ԫʪR�O�w�r�����/�>���)0�ǽ,�S)�cˁ��*:����{K]ryu�q;9� Л���W3Y��i���Y;�P�3�
��WђB�y≩œ��S�]�5C�T,�5+b�巳F���w��$+�1�i�X/�$��U�{����=b�� �׺�>��w�^h�BL]rC'��E��5�48Vg�L�.������h�k���t.�-�i�2����(�X[�U�Ŭ+�B��U�ꨜ���vQ��v!��4��C2R����9X�v/���(n�.BV4�s6*{�e�d�'�S�3Ƣ��������A�2-V��2R}Vs�K{��e��'�B�vC"���u���3�FT�$�e-��YM�5�u�I[�Q{]^�j���:��L��	��X3�d���s55B�{�*���Z�S�W:Œ�Q�7�;.7_��::�uUFV	޽��U~�b��i��^�I1��G�k����eH����woj=������<�*U��ݼ�^��ۄf�<Tu!j��T���=�ќ��ĭ0R��A������ge�c5s9۝�S<�3ѹv(^i��N.���b�����a��ջ���e����)�U\Ea��u z��]��;�s��H[�i���W���M摜�2��jbj�
�ƍ��V����yug;�}���U���lqr�ډ=U��Q�z�tV�;ƋT�-�j�T^���.jj茛=ь\��0�>��4q���3QWBx�{�5n�&oN{��0A���̕��I3.���e�[ڵ��3��4Cv�&� ���9�C�e٠Lֺ����\pqe��{�^<�Qqq\�����{�Wf�ݚ�w���7�5��-m�;1.D��+2py6�k�뺣��{���6��VX���Br7D��[՛�G-p�)�s�ɽ�Y�jN��Qޡ�7���k&�르F�T)��`��3Q�3�d�S���?v���Prs����{^�q����.����� s�*z�bo2�S[�j\���5t�6.�.�N2b��*wrUU[gU��k.��1Y8�5��V����j(5�y|��d��(�%;�&��76@����{~��3�������v5��wWg����YbT�нՎ'Y;���D�ʂ��ޠ�.E�����tL�.��3�*p��v��+Ov�	���y<٬�"�#|�vЇ:1���ԃ�-V���<nL�̘3S=�����鍊4h�w���jv��b����'��,�sh��9}6�_n�!.5fo�Wx����u[D�nX�r�cw�܊Q�G�8������Hl�����$%+4��y�u��Ū9���|����q�ö�_AN�����;nTf�J��-�
��.P���Q�3,�k��zYnl�M���
�^m����O!�����yjl�fo�d5|g�H�r��[�1��9�����=m<�J2$j�h;ԥRث�Q4��c��Sp����=��}�����^l�ڽVst.��Z�9b�M^��9d2'�c��y
�b��j��'��Y�$Κ���U��x;�VV��u��5�/Lm^�eh[��ٍ���qI����ٹ���ZÐ(fdS�{��D�������F�lՑ�",�S��v��yr<�9��]*xE4l4�T�t�E�
&j�f�\��Bm�}��N��j7=���+����9#y���j�V����*2��Z��YWx� f�C'�:2���V=��V�.��1�L3��fo�FԘ�LM���^H�ɣ�p<��.sp�N�b���٬����ڃU�z��##�y����O[���Q���׼�r�����{3nֽ�}T���*�qs[)Ո���_>�{<�*dil�"�n�3�ם�/��d3��iه�s�t�����^��`����&	D��f�s��Ff=ҫ{�8Ș3�&P�����'w��d;��-�L��Ә͵Ӟ%�oqjyٮ2���X�-;��/S���.��6����p.%eQvjv9�ع���}�eɪ����h*��]�}Q��f�n
���s�s���>��3˸�����"xdy;�fpF'�e`��Q�3���Z��:6�
@���1��K4a2�.�8 U���WV�>|'%�3xv�O�bL6�������"�Qg�1o���r�pP�H�h���UѨ�q��V�'pꑐ�����������/'�Xũ�#Ib�ܽMȍ����6�"W*t��\�8�S'�eA����:�:�����é����S�ҷ�R�M+�a<�;�g.E��vu��^�W�Δ����"n4�>�lf����{UWϞ,r�6��v"�%v�٩�JW+�]5�: ���%��C6	�s��.
���0�ިV&UeVT�@S���o���Z��\��7��i�B�'�S��	k�㊕��ڹ��T����
B�Bh��=�L���m�AYgF�r���vîr#�,Ⱥ�sfv-f��ōu�g (�wΉy�J{fv4P������S��P���ܮ��r�a\U��GA8�R�s����P&���q���Xl���\v��k�	��t�ځJ.xl9w-�L^��#��q����ډΨ��A���9�mo1�يqf�)m��c[1����2�]��I�ũ���H�:"t�*�iq�,��y�ڕ�VSͲ{:[e��m��7<!�kճAB���*\�w�#m��ge�)w�J	�jÕM��<=�{}��9�]ѻ�rYتP/�,wp�S=uW)���|�N�W+r�d1�_Kə�\�w,\��'���,[���<�����������/����h_>�B�П�߷+�\T�|o5[��ӹ�~�/�e�]�N^\v�L��<�՞����Uh��Zݾ�������7�Õ��{�ȋ���V���1y�v�GR���.�9�@�IJ`t)0
v��#t�ˎ�<y�[<gL������
B3�o8��Ǒx�^���������tb.�-̬2e�Q8XѼE����o�:�g-$/+��}
b�.W][������$��Z(��pL��kf{�^FKeEf!o�U���N�VO�h��T
bw���m�6�8 �ٜ����잃s�d�T�P�d�{nE"�aiuF�[���K:�]�s3TX����7]���2r޶K��aސL�T�C��U�5�H�Y	��U6&PƯ�-�ԧ1jUD\�M�M�W�ԑ/.
��o�l�}����Sl	C�35`�3�롇��9#H��;�7��`�6�	�3j¡Y��%#�Y�C�Gf�6���\�B넧,tk�癦A���~p�"���9�\m<3�v�8�ͪB������R��٘yF;S����������8)x��\Ť)����&�o�>T_#w����B��V/t��ĥ����t,���·3e]��Qq�'����e	�o�@��X�;�N���ll1q�2z0@�*�z���;њ"�ԃ{��A�a&�s�	]��v�3&�mٸئ�h��3f.A	�i��(_o%�Wd�\mF��4�M%����u�O'�����r
*.�㙪0�����1[0�u4k����7�wn��	Tm9�y�����H9�a���'0�MmT^L.5`�^�3��*� ����N�+��)ܾ=�д��_*�뭎�k9wa���˒w6-���]��e��UB�[��o��rκ`���#T���S�X��W�' u��8�:Me�u��3�-0�H�rp�{�\��T�}�C,﷌���w���a���w�Rjnp�&r��\VO���dsGK�wSf��S���S�� �1�u��2Ⴢ־���jt�TS�WcdmXR�,��5i���4Ӳb�9�����.�i�sF�<Z-%@㽱��H�ʱ����M�q�z;��S�vޭ�c5��Lӭ1O&�u63/�]K�W}v@�w{n�(M��;y}�O[�f1��	����S���r6}���}���Y�2�_�'Y�i����r{��6����
î���ʡ8)��j��ǂ0����˸���y���T����8�7\�p�o�l��\<z����kn�gf� g���Õ��S�9J��\�(��Y�GZ�}k5�N�Q���$Obn�p�2�ɇ{`q�WWUWu;p&��'z��=<D�����]i���Oz�X�P�WW}}*��s1�
ȗ���� �MM�K��6�� w*�RႪ���T���P�-��w#Ǧ������].�Ψv�h؀C6��t��%��U�L�+2|{�m]m���/0��B��T=�N�����OJ���M�Ѭo	rQ9#����1G31fF�����x��m٠'�-�4�rZ5�μ�w�YT�3uN*6Hp��Zgm�d�]ϯ���U���q�^d=�+p���w_e��c��SÓ��aӌ��N�i����i�E��y���;��m4���۸����pj�^I�L�#(E=nLoS����i,=f�-o�]W�C#���#z4f�e�t3�Li76b��f�]��&/1�e7+%���ky�F�30M����IPYՊ��Ut��f��Sԩ*�Pow��"�X������� ��e,'���^�5c���9��«��,FD��t��O�Wڦ��M=������țݍ���l�MQ��s�s;v��n���#�\d�7�(�K Fݬ�˕%�4�jNM��[f��k��\��{쌿9Bܙ�ۙ����+��Cvg3�6��3<��n�4	���r�;	aI�V�=/L5�*����vb�:Vj�3�;w�(v�t�[��Π����=.����(v6�M�kc�ڣ�3f�5;O.��-jvz�-�s��w+���I���aٓ[�˷a�)\��aƭ[���Ȇ&�A��vfC�zW�Y.�t'/���ʉ˶��:�)u��Y������[�.�:�����5D��oM`��v�9iރ=S�՝O*�Q�ڦ���B#\S�T���]Nj��d��&D9(�@�^�f�ظ`���4,�7�ol�L�ۍUSI�hAZ��ν���{�o�A2�շ��CQ��`��M&t/p�Ŋ��Wf�>t>���D�$/��\ʎsv�vGAJ�9�3����Q�`3X"/pKA��Q�FNvMT�Q9$�£�j��#[�����٩ڃ&v�&�U��C)9�{8��������͊#V�[U�9*(J�jw�
��ٱ@P�"�j��Z�UgE��K5OFdM�$Z(H�.l��ZG|Uι�"�qb�m$й[4R��e�2��4���e�,�����p�y�L�znPǌh����q8�v啣��%c������;�L�7�
�7/��jiup�1��z�W�7K�6ؙؗ�K)M�v��㙜*�ݓ�j�U�����/U��.+�O���q�*z��K>���qnEy#z�F:&@hQ=���:��h����f��kv�/̥}�9���ve�>l+ۑ�|ԋ���V���t�1���O2D;��Ӫ'���s=��3ۯv{�I�qNꢯ�j*;q
��ъ�puun��.9M�]P�I9Q��ܘ�ഃ�E�ɽ���gr;2��Ր��O2�U�Wf\l7cS2��=K�H�c�st�uc2�8�&��l^�e���y�5�`��������k.����V�V�3P �ҁ�(,�ѝ;�;0J�᧔�̗�	�Do5{��dc)ud��ʎ�v�{oU�*��y�hțYUtm�;�1�`��gT)k�Q���� ���!%��\�P�����G��|�8
*y�zV�]ݲ:v��<���T��b���H����YJanӛ����䭗�Y������"��Y�O�Cl��Q���Z�B��S%7S�� &�Z�*��S{#r#3n-���9S�����p�! ������ǵ=N�Y��zcdE��ڋ�Uy���"+�٭t�ξ:nvTn��v�f�L�z#F
p�|��\9"T�U���T3�K(�;��]9��Ը�tPX�k��w+�"�g����]ubq��o i'�K�ސtp܍k"U��H�\���\�gd8�'�V� �lL�\Vb����F���A�U����ӗ;�@��@��6��U�K^#��\�N��*��i_G���8�Ú��s�1~U��ضd��.r�uL�lr�|[
*�jd�x<ha��d�m,�u���:�4E�lnt �ƛʒ�ꆪ��b ��n@\굤�t��Q�����z&f��ޝ&��wMʘq�Md9"p��f�Dʑ�Ds��u9����݌�vzݩ���2z	}k6�si�c\������{0;���<w�����s}�>���3L�ٽ-J���V��+��'���f4eC����fF�8mk�\����G#P�wf8���f�9{�1�5�
��E:4nT3U�s�v�.�e[v�
���P')l�ě���bv�TB֕^PΔ��2��p+�m0�T�x��vh���k��/S�v����0�ƛ<��rnh��mr�6���|�e���Yaf��s�h�S1�K�f��w�%�59����t����AmnPN�Pf�]w\�����wb�f6�(��ޅVm�5ݹ�c f�k��V�Fꡮ��ǉ׈�&�6�wtڎ6�؆F��p�w$�xe�W�l]dK��"0����BD�KH���q������q!a٫�p�l������/a�Y��V��U��M+�q�-�\��ph��s!����oD�ѕ1|ͮ[!m/6�=����%E����꾋�7�USU�Ô��=���e\�	u�-
r^ړ������N .X�;m�=j��,jyt�Wo��Os�wZ�w@�� �h�w�-���%gF<sB�uE�ґ���22��Prgh&� әR��F<����Gl��+Y��~��|}7J�g����W8�d�n�H\U<f�Q�R�ދ&�!�b�G��Iѳ��O}%�m��zEκ*�M�zuTʾ��fb��^���݊U��\���S�����U��k����&�t�'1���:�Յ�6����V��3�L�L,b#;$�M�_;����]�c�1��u͵$���y0�v�D�>�
ә
'Mtw*�zH��j�������� N-b�Sx�X��J��bEu>��L��hF:h�YGl�*V[ìS�pT�tݛ����}Է���sQ��]׭ޞhߴ�CI�g��I{<td�8&=pu�E��.�l�ގ@>p��{2�J@�wKnI�#`�;5.4�m�"-�у6��2{�{ۍ3&�c7��͚�Q5�k�U���W_y�m�[�v�\#3�5廽���(��)���xq��E�*��&nȘW�{�E��8o;Y�ُM�d��L�L�勚'v�Jȱ�4�*U�����)EM������6WE��T�����N�î��P��º�;�2N\�\f3�]qr�����*pV&�V6�0�w5�R���񼝃��F*�f��F��t�v];#g&(l�.Dv�T��=.Tb�3Q�󖺪��8�`��3n�ڗ����)Q����H_NByܰ軱���H�vE�A�1jrg(\T�0�jz�oL������J�
낤>ɽ�,��\��i	��;�~��Qǅg�9꽹��2f��Y}�7��6����'�έt���<����x�������P��(����4�T�1wW���'3p�Nw?f͓[d"��w/j�n�mR�LK{4.��}B24���8��l��6�XN2�{\�t�"-�ܭ݂���N���D虡�{��՗t��U�N��3��f����i:g���n-����xut���9�'}�F*5�i�u���O.�ER7�U�M0!�G;ou^��<J����a��gp��Fs�Q��ޞJV��R}y�ٷSU5�b�S�-]�,�s��ca;5h��x����F^��^l�s�#5ew�����v�Yqջ���$Z
c��O�v(����ĸ�k�*�wUnTʎ��`Lp�K{c��w5с�*v��:���T�^��Cwl(��V��yqق���r#f:��	�Z���77�Q̛{y4X;�a��y�%�D��^^��P�SO'	�͝�yD�P*d=��d��̕R��@��D}�4�h��%q�yw'�[�D�����R��y�gi�����qx0�yqG��|'m='b��Gz��ǜ�
p65��������r��;�l�9^��{��)�w����qp�m-�
.�1yDۛ�zՌ�R��jM���EGF�D�0#~c;�����DEՆb5�eWaN��#U��&^F`���	\ŝ�1"h�����Zzݨ��LX�N�P�Q{��XEß6����plgJc(r���^TU�l:ջ��T\:�ʝ��p���Z�ҙDF<B/IF�Nx�6��s1���[�7��,S`>l���%BT�6�V`M��yh]�#�eV;�6L�e*��v�n�������X��=4��Ȝ@-�d���;;�+�3���a����0�:���ϴ�h�� �I�$����Nu���t�
�dH��+�����s��0"��pL��Bp!��YUN�Q�6�e��W�;ݣt:K���.�.f���bU�5�E��
��Omڍ�-QfiT[\E$�t5�2'o0�-��[�l��%���6n2����f��&��f���()�ζ��5�X�Ș}p�.���U8����	̑��e�G���G��B��i�4�	�d۩0r֖ظ�y����fs�w�2�dv�Q�ח4��ïrL��~�W�����ݨ���v����]Vt�_9��^��vC�ewׂbﷻ�3a>�<��F�p8Ǖ;@t���if:��w]3�n^c��U�'�^�V`{}��\=�{�3�wg�ۗ.�v�[I��d���u�=�r�i��k�vɌ=]����;*pw�Q�35X�:31��x3S^j�D���ӵ����Q�}]a����q�@J詢�њ���j�7��{"�ER��9!�K��$t�F��+�[�F�"b�o6)�F�^�H��:3�v.u�<�Dmn�tk�L�S����u8n�I�S�]�8T����g���ݶ"�����2̚�ۻ�qgv��ص�`>+��޵'.p�9}&����5�CU@=�=y�pi<��v��6��v#�wgd�ZV�1���
��4��*%A��xgP��;A�b��[�U�7ζ����ikʅu:�&j�恊1pʽ�u�&+�I�q��%	�{�n�^�'�[F�n�Uqn�g-��Vk��B:+|9�����d+��e���`�8ep�%�1*�Z�s�;K�5��Pna-ª�vfa�T�W3]�:�3��#$v�#��B���9C&r6⦭'-�i���3���2��;��������9�t.�%uj%��Y^��wj�����Z$R{=SE�z�ߗl8�K�E�I5�=�;���v��RGi�]*s�m�b��%� ��e��\�j��p�{i�ٚj�؃�&ɭ��s�ssZ��k1v�3m��;��\kv�j����xA��[E�	u[[��Np7�no%Љ�9��%+X�qh��}��{�Lɻa�)�T�H�Obuf`0:���bV.��[��f%�.�2f�99�ۻ�ÑS]����͞����2\H��dLUr:��r����f��h���E��^��J��{ػ�*V��ƞv'&:�V����8f�yX�������g0\"i�2d)���t�����KR���xi{��,Z�&�oH���o� 7o�/p�Z(M�b�#0��9�����Rnz��9Kds|1hs=ɡV��sHɇd�,|���D�{#����ZP��,]mU&��b�6�E����3����
'�^��3�]uf�U�U<s7ۓ�9��aH'T]�dU�-��ٽ�;LY<��^byv���X6-;��Q�kV��t�'.u������'�~�����^,у�eJ����2\�bz.�U_q�J�ы���Yg�X��ث�w�eu�N�VV5��Xȫv������w�)��ڍ�wq���D�6� ���۵c��V�N5{=yՐݖ��ɾ�9i�ʺ�Y[M�,�$ܮ\��W�8�ʵE�U����*�nL��α�U��Ok	ۧ�VcvZ�~��)�Y	yD ����"�2# �@���lcX�Q�+sV5DF�F�m]+�*),i"H\�Eܫ�h����n���k\��ch�L"�sm�\�lV�qάj�Y(�ZeңQU�Q�E��2kXMITZ�����w���ǜ���9z��r��x.��å�c��~�M��>[Oc�~�>��5������&��w�����L��]"�����9��K�?�"���_�T��-.���cw���1_���ER�8z}� Jd�t_E�9�8{A��'?���"LI+t6�s3���I��!W��E�!�S�jb����^�xW+z��)uP��yc��E�o���u�ϥs/d���DW�%.kd;�$�_��}^��.��d}�������x]u���yE�������U��Ot�<��[e���b�H�yv�wز���G��� ���d����D�H�Mߛw#��_]j��Ow�o:[��>�w|9����|���!�8��26j����s|t�dqjh�r�\}9Ӵ��ѫf��Vȍ��a����tcݝ�wu��uf�b喻�T��6�9�ޕ,�xw<��2�A��P	̓�Xt���:ڮ ��N�R��ܐm����4bG_]
����+�I}��#�%bw������H��J��q�XSd2-i�mm�xc�A�ߦv��7�B�q��~&lEL��Yw<D��Բ����$��A����d¸;�6�]���4`�A��{D�U)��r��H��2u8M!µfi)�6A�N���Ty옵���j�*]��o�ˈ�ɟJ�~��3LC�<��㭵:�ށa'�^��ӫ&]�s�fR�Ur��e��-�	Q^�^#&���,��������u����$�̖��=|���j朎�ؓל��t�����5c��e;�O)Z�E60�E��ǟ��i�jr=��Z{-�mL��9]��T�x����<^�hZ�p��u�̺�ͱm�������U>��2r�}uʵQ�n�)�N��۝���%�@w��'�1��s)�d�9i�r�d���{�De#�g�;�'x�U4�u2��>gS��ڼB{m	v��Nԍz���CE"�.�yA���_V �<^���� ~���ݢ��k�c�J(��q�s��#��{�ƫP��F�[��VX�b���)�� d��_��7jV%W�R7a�.����\Q��pa�?���<Mm�^IkƝ�!��ߏ9[m��9�d+���ʵqaX�M�I���e�P.��`z�=���M��RMb�
i��8u��� XO9M��]h�9���}yK��p��u�I0��a��:g{.���!��te�y�Q��l�{u������Q8�;e��[�
�E�8�5;ҏ&�j��6oF�5/+"����Y�wR�wAQ� Fhm�uu�����K�cf����� �+�&J���oș?=w=jP`Yr1A:�+
�D�z�I�զ�1������2�}#�1��;
i�_TZ^N��v��^�����(�=#F8��>z��������v���̲��lW����&�͟Ff���3[>�^�򏪽9v�r���sĲ���'|p��e��1l���V������hbHx��\lwQ���w�����u'���*��Z3]�]4IF����0l&�ӿ&]��3�J��4z�uFE�+ڳ:i�ή�2�z�,o63�:�<��C��� ����z��96=P�ʄ�M����4�$sf�tu��8ָwV��g���.�r�6e� �"L35�L&
HQ��k�U��ѕ$	C?��.�7"<�a(s�"��{�^�90�fK.h����F�샘\�;�D7`�<O�O;�kkAM�3��K�~�T�=����D���\U�*�+��.v�e�+?Z�^6�H�C�����3�׸K���b�� ����RT���}A�o�{'��(4/w�����W��H�m��9��6�WFryH伴=^�n�^��"Q]�z\O,���_lv�;t����P��i=Z���4w,tz3\$�2���8ܻ���l�� ��Pv�A%�E��O{F�&��v�GV��`�oݧ�!Vx�R�Ώ�R�_-3Ѻ]�h)����~}�� =���+�� ���?�����{������	?�%��G�7�T�B�뎺�5�x;b�?k�ӿ��0���)Lx����"k)�V��w�/��kk�6��ژ������C��éqx�2�9hv��׬�1�p�Lc�T�/�u�B��k�^�&a	G1��R�B�(!�P���s|�;��_��-�I����x8�J���r�+oo�^)}��w���b|��÷>��P��^#H{w���*��n;�ԡ���&���o:%�y��꾡��o�ۦ�]�ש{O��gXNыV��Mn����ڸ�-� �Qs�K}�[�;;<�������v��)C6�M�_�{<�xZ�*B,�.oߞ�ـ�������⑃m���Lu�,牬�١�sH�/YJ�;*G�z�<R�z���S��o@�w�!mz��8�ש���H�;��(���޻��U�ٯ��Ք\����џ�@� @وP�� Ȓ*S�{������NO��[r��~��?����b�l�FAR �-�;�E��]���~C����9"t�?w�R4_}�ų��|���{�|/�7�m7����!vW��ľd_�|mg��}����ɐ�w�P�̲?����]�.o�~�}������?�i��Ś%p���l�p	�k��?4t�'Dܙ��7�='�9X�����_C�"�J�_E|��x~���P�ӹ?���ig2�)���gj,^G�{)�yx��t��@��� =��Ǻ
k+.�����_r��4iP@>�{�Q�o�֦��2������L ����!��w��4n0�3�b�uS+�V��9���!���.��<T-�5b�(yQ�8���ba�� ������B��HR%I3���E���V<�Z���t�Q/a�v��{�/�۴��z�A6��&��Z��Z��T����E�z���-�+N�Q�T��I���)����j0u(p�������5mN�2�|"׶*5� %��!�9�og $3mϹ�9��{<{l�H㯠��Tt�=�����������5��E9ұ5��l��d:'|^<��x*��ޔ!�ͯ],g�N����mi��3'�`��mO�S)��/~�о~��360w���үӦ�%9Ny�E*�L�|�
���ٲ��U�6��7���S~���N��ػ��g�e��O�;ѽ=�����٧�j
�h��n�iȲu���Fr;M[y.���u�ɻ�Z�A���/�q�:f<�}�&1hn�)ʜ֍T{b��z6:'���d��U��c���
����GݽOҧ9����O%�fjӇ�ks|��+O�<���_t|���K+��A����	�<�p�N[������b����3�Tj��;����q�?�QS�,X��f�f�r����z5N�OoJ9�*���kU��]wk�]�^�;wu���(��8n�}�'/&�/W�]��{�v�#.eg���	��lx���k�;����Ͽ�?#LU0Yݑv�憹��������=�gUyc�\���8+DHWb���z��=�8�fl���o����$L��G3�eܶ9��)�\���uZ�-IY�w��Ӹ�;3:,�
�o9�2�_q�Ggn�rW�	"�X�Rnۮ5鳕V:��e��ˡQI���zr�@����{�.�����X�nN�l�QL�/�|���S���X��B�<#:KD[|\%�|D#�yN��uK�l�ҙ43<dU$yOF!�s|���u&>�y.�k(��ǔ���|t<�3�Ѭ�x���q;'����ew�v\:y��P6z9l�&6�s~i�u%3	�Fx>��~]kȬ��By�N��T^\��&"�e�X��F6Q�"w
�e�O�,�U�ጀ��_��+�]@���:,����PU���*�4r��hH�9�$�EՃ�F�։���e�MY3Ҁ��(��v�*J������Gwā�e�D��Z&�4���OO�}6��5�![��+��UE/^eQIΓݼ�F��ވ3��,�pۑ��3�
Q��e�ub�A'��*h�ӯtO)���!(S�Q����4>n���%~M؆3z�t�,��+a����y�D9){C���7O�g������~�[���[�%�ee{뽔�_�ӝ�j- �}�cQ�c5$����DM�R�/h�����o���ޛ��AHv�
2;p?�PC�~z���_=��ΤHb��ĠC3H��|C�;��=ĵ�/!��������*��J>����\�,N��a�����X�jٱ:ZhW>F'5�)�jU����G��Τ-�޿�S<�H�p	�C��_�t�v	��''��K9*��i��8�+��+*)I�F�y�sE����˲☇u��eO,������C�̊�!����3cm��`�(;�3�S<�$/�Ri;��T.PyIl�=��u\ad�-۟�w���Գg�ꁗDX��"뀇��Mx�!##�GK[B�EdYZV2��tP)V�2-��$��� =��O�y�~?���/���#���wx���o���5���q��CyG�v�M�߻�O�'���a�G�����":3��p��ضsv�E��6lwٚn��8mƫx���XB�PY�Š�3iC��]%ٶ���5�V����7�+#z���b���P�Ti���u�a�f_��{:������g�L���]2ڏZ��<u��Vֺxj�;bv"��j��U��7Xu����6��Cp�E�cS����h[h��ʰ��U�O�Ba�ԯW��Uzg�R؈G���v�zsag���1a��E9]J�"��c�ⵓ�!�.�4�|ۼ_
��ݞ6�Me �ƽ�B�;뼘�Ve�7^�j��ݖuW[-�W���W�K�m��;C��&�q��D�h�Z���{sY���v��kRfŞ]sN?�  @* ABPY �'�🯼��Y����4T]"t
DD����J��HB$��$$�I$!	)^�M��[�����_�Ϝ}}�,���S�ŵ����lc�ċȼ؊�E^,x�i	�h�dV�ĭM��37�͆���5���x{g{�s��#��Z\^��-S����8�V4ujɫ�Sn&���h�<W�F���fx�J�a�@�"�Z��f���N�P�(�m�[/6�7V����Mg�l/C���m��T.�!=�՝8�N9l�1+�|�d���6�W8��j,T*�>�����3���eY��ڌi=�f�ڏKn�4�}�!�K�D��/P��Æ�1��Y��Љ��/�hݪg!��k�NWlZS��HfN���8�`�Z�G.����DDw����t������/����w��ʙ�0_3� R�E�`�"�b	`)b!`� �*� !��Ϣ;7�x�	*���>+�+W������Qc������@a$_�B�������?޹�f{q��k�z�ߟpg|��]��H�����������\��`e��$ӔeJPV6�5�\g9���r��i!�fm�d;bX����/\�y����EUk�|���e�p��>�w���r&��}���W�����⾑R������ߙ��P�%�Uhv�dĝ����ߏ��9HN�Y���i�N�X�*V9F$�$"�
@�Cc��˺~���幝���?�j���Hb,P�o='ׁ9*�IJeWI�Y4��E��+J'dk��E�4w:���^QR�T�i��I�AZ�R*ގ��Y����e>�x+�pI����s�'8&��Sy�`�� A�0�Pd�[k���Q�dq�0"b�:�b������g˥����#�y~*��~��t^���oϝA "���'������&�o~M�=�^��Ӽ���9'J?o�?<'Sk��|q>;�������i9�Ma1�M>-��au].��[	.� �'���AɅ��7�������)RK!R�G�Pn�N�Ѕ0�,)z����`�fcЦ�n�0h#��{����Q�����#%�F�B�����V�E��f(/"���2���E�nK&�\	ŕB��O��P���qi�RA �]f�3d�i��Ų�*�k�V2 ��`���AJ���`�E.$��;]?�⺥,��P���ӣ7vRY`D����H,	¨R��A 2I�ZlC�m5��X8 ̕Pm7j9�6�H+�-z\8q��"�E���I��=Q��ʴU�*�<햭��\Y�`��	���]��'$M٤6\�taBD�n��� '��h	eR낎����dڼ�Dw]2�Z��+
ޡ�Ix���
C�Z	:I�m�v�o%��2�1I�����6���5�%A`�/����1��o ���`4Ur�6L-H��Y=B�9\��m���$b*�n7 ��pXMU�ݗ]+@�U\ћ�p�
D�4�W`֌�!��l.ad�)Y
�fD�L`�&H%���y�g������aW�>`�y�FQ�fA�(���>���z)�.��E�`�1��~���ٿ�Lti#�c�i��s�� �5ԯ,LE����.G��O�f �]h�H&q�C;���29TP@$'��3'�����
kF��V$�c����02�{s^�RYpZ�_E��3(X�21uPUT�C'�a0g+%��|�n^ ���ɘ��Xna��u�6��W��p\�,R1�U3q9)�"׋O@��h�Y�Y��(;g0r�����ej�׃�ĉ>�a ؏���
�;�e
�/%� 3-�Z����r̳M��?�=���xj`� w�l��Č�Bd{LKy�w�Pr�X�^MW��7f-Mc�=�c��+50VCi]�U"�k�I;���l}�0��Ѷj:#�aV�:-�!� Hk��#�w��+!aI(A�w\��#�'�9�dq�͘�E���l�
DT������vX���1��ǊD���l�����*q<\Ga�$0A"��*	��X�m�*�Ͼ�
�+��t���3�	��-j���NձI��*�㻘=�(!EE�{������AX�E{�_4�Uq���*W>��0R?F�x��j_h^X���}[v��Di�e���<q�i6|�L�(C�Q]�$�j%Z͑���
�������I��e��#5�t�P��ZQ� �HV�j����p�� ���&�C��'r�Nj��Zd"汰 *�AÕl�A�#��F3��!hs��>��@��H�Z�J�Oe�U�>wS��-�w�a)�C<j�ţ��0��8��C&�)��WV�O0��l��U[p|�'X��������� �n]5��M:�0�� T��f"�Ij��Z�t�&'�3
qU�'<'"*	�.�;*���SɄ�b2����m����U5��F���B�&�X(06VR���ق�YX����sy��-b3�̡��誊���F�I�S�5��<��R
Cܵ��ھ��UL��!Y�λLR����톙M�(^��m{DY�(�P�(r 	T��O{�
f�CA
���N�L*n:��H� ���s|/J�e0P��q�W7���n 0�Pj�Y۰-�;(�ϝ�i箧=�J��t�<Ic�;�:�0�aX坉-�[w��PP��8��Ҷ�K��h��$��<�Ȼ�K�6RJ����>s����͵�{hE�Tq���0��a�b �wTe9@,m
Y�=�0�Q1N��q�D�9U\���Ӎ�A��λQ�U`���If��!)J�%�
���E�^3�T�NKEq1a�A&|�����C�%C�V)���*�q��
m���0f"�#g�P�U{.��|����а]Cw^Þ��������f�p�����A-���-�6�F��v�a�g�\Ĉ&.����b"�/9�˻	�u�ı=N2�q��c�����<Xn��;q�vߒ��G��߈;�H;لc�ǯ�[�hW���u��uۅ���MB��*����Eڅ�o���6Ґ�Ë�eђ��x�^%��Lv(�{� ��2g
V�vsmܪ�O�v|S�^�\C7�a�J�l�q�[4�P�I���AH!r.��&�,���d�Y������V�*�,˽�M��x6�1ʋg�+aX�Y�.p�YՂ��K������ �0u���ʱ��}-�Af,�$5�*���,A*J�ܶ<JL�n�ɖ���g+=�q��F�#��e�|���&��w^z��.Sr���&�2��}����Euwlj �����s��$g��@@�T� ��7��Du�����}���QH:|��CF-f��c�%�;D���n��Vu*�/ȩ�$�>�,mT�Ug���:��7��^���U_<����(�+����]��D����'@�-�
{J�`C�e>�G^H�Dä$˅VRO�T2:��u�aJ�,�dܛɢI�w���9�'��=��ZVb�W����$v�\`��PH>��Q��j��9�Wx�L�̱8�-���Je3�	\�oĤ"d�]�A�>2���(ke�
BB�TA�Yj�<&t���شzL���gx��C���h����R��p!��{��2����ֺf�n� $<ʝ��q|��,��rT�39ƃ,{5�J����ui�7�&�]��%��ȳ*���Q���0�#pZD]IR3�Gt�\�(�"n[hH�1�a����^�K�p�ƻ�Uj7����-�A���r�ļ;ڡ6Z&��\�ҹ����~���+���gT��7{��ݔo���k��X(�CT�J40pis]�#�5�����U6#���N��y��,���l
�a��B��ק{� ��A��e'�h�c# p�-��!�ɡ��R���5/�����0}�1�bHK�M�9`��Gi*0���^��B��g��-�D-�L���� -��H��K�Ƙ�4G��&�z�/m����h����\�囡<,���]ȱ%�R$��DD�i�M�UXR+2(U�7-�7:�$�c�P)..�"�F֩[P���� �|lH��~�D؍��g��v�K�[�����!IU�,���(��̂׹S��N=��#X�q�x3�ȉ`��\܁��AQai�0��\� �f/wʜ(�S傠=j��{�]�)wR�b�`����V�c�iL^�D*�]�	������w��Ҏ3 �c*A!�]�ĞK3G��%��Eɋ��!�\\ar���9�@��>0*��ڸ���8(8�>�+ѹ.�W���ֱ*���ǐ�X\=�C�u(��T\�ձ'(�~�9��K<�= \R�b=���'(7bB	����	��c���Jd���X�r�,��U�9�YQ"�j"�E�)2�*f	15)X�H� B�cq�)�Y���*.`T��f��F]��*/r��-���+��"6�/��p�`̋�;܂��H��Hwf�x.��$vId��tUJ��
KCh�8)�3W~�l1�I�oG ��3h]^���<s�� %;�Z�@���ǭhWc�>�6����𠜭�{ສ&K�j���d���e8��S{�F��~<C($t������:�SLD�/I�*AW)I��.�$��a�P��:�/�&�Ɨ��1�F)����~6*RTR�$���MW����*�%���8]��[���Ĉ�J�L�tn��ػ�T��-�a^x�b�arE�ˆU��:5���y�*�e�&{,vU[��81�J=�|ҥ:T�`tVv�6Nݷ)�|�*E�5���
�a$Wj�`.��':��UI�a���%�&�!�V#��J&�J�E�%LL5�D�(���w5�ɟ��:kD(؅(��Lje�Ę�qᯠi@�B��U$�aT{c�|#��B��b[U(ޕ^H�'` E6��e�h��"�gc����S$X���`�(�0k5�I��,ƨA��Z�E�X"�έ��7)1��dNH9P�"!��%wq��\X��d�%.ȩ~�P.V��,l\��P�#a* �iXUčޕ���X�m���r02�g�����"��`Y�Y�՞m%`H �g[?�`5g�8OF��&(�z=6

�r�n615n�i���Y��T`�1 �{A������dd�S��r5J�\1#Q9�h��%P�q�zfj�*��H`���bK`ff���J���6��"��9̖�0�-Ӽ�k�
I����heY��.PZ�a/��I#
���q��*�-:e���J�#�5��E��;�!.#��9�T�T�Ww�i�:��TS\j�[�Uk<	w��,�\�C�
0f�P榀Ѧ���J��5��)�07�<��e	r�YT9�H`ź�>r�#%�\�z|
�c&)J.�$��E�8Q�^��E��
�Ҡ�(�&��X�_xh�<�M6��AA*��Ѐ11-H�$H�oA�*+Ʌ�m#��
���+[U�=���X2�0m[���T"���FT�ن�7��)L`�UP�,N�s(y���6�7PˇU�6&�_o
"+�I$���9�
BR��F@1&dV��Hğ!���8]2`F�Z�j)���t�r,A�������
DZjĒ,R/Q����"0i���t
��%�N����2�e���l�GBc�<2�(�>�0@�0�Q�8aC5&�(Q�d�j��8B�w�bb�\"kuT"�2��2tއ �$��{R�("lLT�Ia��3PI%�� I`(���w^�N,��H�-����U�a�F�$�Z�-��3�8	W�ԗE ��m gd��E�X��f����"�B�V���c[ѲL2��bB$<�����-V�,6l��n�U ��`m}�`L��
E�D��{�B�6�j�h>(࣐��Q1ch�&Q��B$Bv.��)��
������A)�5���H:���(�p��/���rȫ��L!�׵��|۹�bv{ �Wa�m�� ��TY@N�vq�/X�v畹��j�'�P)aDn���U]Em�y%�;aP\�� K�S�ҹ4�CuD
QYŬ���A���"�T��aPA(���q@�d"�P4QYu����k�&JYpCUH!&Ӷ�� �ÿ�`�v�&'�ݣ�����8�P�mX7�����uO�|��C�ta~<,������xU��i@ñ��k��a[��5�j��to*�
��jh��[9�a�cS�{��ʊ6ՠ��+]Q����l@�֥=ߵ���T}20����1�c2�]�.Gw'DS���BDn�������a��^N��Q�
��r2C�pD� �(�H�wڒ�:�#��T�����KI�h�m��a�Z����y�ţ���[�:4���~BC��[�a���P1�Ygf������((�b:g��! d�MFv���1�N���(�$�8�D-"P�v�隖=��7'B���l��*hG
H ��۱7;{wT�<s�m�)����)2��#	*��ŊR$���sC^��թ��;ٰFŁ@���$���)2�
X�(-HVM�@L��v24�(�i�'hl;`W�W��ܡ�H� �(��3P45.��&����7�@$�D�L��<��:.�$���Th4�F6y�
v(��w� �`�i� ��Gd� ���м$�G-XBP)@l���#�V~* ܁��1=�Z�I.$�O:�m��@c���1%UANX׳p�*�]\U�`�T����ҍ�Ѓ}u�;U6#�(�$7 )@�C�J�"pB[T��0�V�<9(Hs%6C�Bg2JI_vs�n�o hB�����2�Ds���T�jl����p��<�AV��A�%4R�j��v&�cqbl�6 ���H���M��tAC�>�&�H���b��f��Ň��N]-�.�>(�B�86jX�3*��
i\
��XN�Y���pE�l���Pp�9����(0ᕮH!�f
ATT��፬�������P)NN�緫�"�M��F��Ñ�ㆅ'���RʠY31��wA�HT�NH)�"�ŋ�"@��p	 8e��d�-�+X� �R�Ef^*�!��dk�n@�T�T`��
E�J�Յ�+*L�":�	>��bpK����b��7��bª\��M�y�M�T>{:U|8�Ǩ(�Ć�g�AI�`�0��J�����j�r�Tsg�l&`�!b��kY�0.�7uReRL�TC�P@nOy�Pȃ+W�@�:����) �udV��d��(m�lh�Eª �k��ӫ��I�P"�Y��Q�c�% T���tR&�0�iG��%�@���b'���V����$��P³,������&�^@����' ���S�) ��km쇛�Lj�dQ:2�HSFP6jM�C{�##EZ��ђ�a��W�L��y�r�*�B�Ũ
�N�8��kB*4E��TtX��a�4��k���K<�'�����Ј�UTw;r�Fvn���e�q��'�hB�XE:\
L�x����cs���`���X�n����F�`��ffe.��k���GP�wi@��έW��Y�S��_F�O�8�.A$��0bM"���i��X0!�D��Ӽ�1H;R�ݖ�C�{4'F�ss���YU3��mx �̘6'{m�r��/ֵ��E�N���]v8,�ɔ9�m�9*U�q���TC1�Web���fF�ɓ���Ԧ(�����F�g��0f�Բ�e@��bS��qA5��]D�� F%��m�2���ɝ��T�T2�°(Yd+�+�#�܎k웳r�Na�0p�B�u�����~�j�U�U�i�
�v����O�}�_&�&�]�A(P�T>$�
ɓ�G��
���o]I���&�e�ɮ�2���>��H}>%>����p�q	��"��YKxZ��d�6��6
U������.��[V�����
xf&g$��G�F�E��BY�DTA֎�B��^ږ7vR�.Yp�Wv�#�V[� �Ys�`�'*��A�M��`�e_E�!�W�����d�`�N�8RLʘ�#�[E��mlЇ
)U�!HPlTPiaff�ф�T���=��-x�j�*�g��pgj]`�}���ə�scW�$�PxW�~��Vi�ʅ�;�`c�4 �W��wV�ˉ@,6"X0��VhK�f ��ɝ�`��Y�!ɔٔ��R#�V�Bg�4�*�D)U
0r�T>�~��EK�]:���ŉ%��BJ�!��ݶHR�"RH�v`���h_���k\̰��[iT���|�&]�x)oM:mR�`�=�UWR��c�⸽)b�eT�����׷��̰�܌��F
�xvy��F������mЈ�5�*W� 6+H�U(82�}0���m+H��V,�zHCk ZVB	��V����5
�wR1gfjNe���rcL42��|B׋e�u�3�Pvf)E[�Ȕ�Z[���Y��;��b�n�t��)��i���;���^
�R!�$t�=l�c��g$ol2��umi�nit{��4��c��;��4{�Q׫�ޔe��4W-�,��~fF��BeO�Y7�2`?�<�T�KP�ʠ��jqf-���h���I�0�}�H-�mH�}*!%]�������A�	6��8m��2E�R@��A�R��Z�V�)]��!*��V�0h�B0�UW�L^bu�{sT�$�W�%�%Jc�<4�S�J�&$��6 du1��DE}D�OK������A�#�c��B�(���0�Ǫ�B�a��2�+%Z֑�\�ˊN:��y�d��H�Ie%�A���ȴw�����V`�FF�7&@��/������+g�w9]���n۔�ǿYު�F�t�i�0�e�籕#����a�[�^��#Y]H\�,���l�-��q�)�(�'Oژ&�$[��(�'8���jӍ��
��!kR�dI�	u�(1��+���|��*aWrࠍ�:�";}�[�#�;(a��{�0�1QVE�V�R �vQkj����fĒ^���Z�d�i>^mK��Z��CG�.Ś
�pT���R����?�X�ՄI�D�R<:���(h��y.�S���i[X�N�r�U���b#j^���\}3����W��b�q�C7c��L�N��A�e����'U\�g�(0#�i���������zRp�R�@�k��s,������R��6j���Ɇ���W���p�v��N��I�x�V�e8Y�W�<]�"�-��mXr���7�+J�c�!%����Ɏ[���E&�Ε2T���H�i:�X��wJ�C�w����~�����Ӝi�}&�X� �Z�4�⣖e"�#��C5e��
`;�gd���q-��Z
�]ĹE#���3�%x�`g�F"���D� f[��ˣ�JXIK�t��I��
α2 V�E�����۳_&m�] ]�Yb��q�d4yֹ�O|�*�Fӎ��:
ĕa1��
�-��^2t��)B�Q���䛋oN�q�1f7��0��'Nu�{h��6��3��S%�(ê����E3���j9xl%��"#����̂.� nT��<-�/*l��*2� e��b`��lؿ2�x��F}�u��m�穨R]�U'-O�%�w�6gr�����F��n1��܂��Sf�GV��UW�+�+w��R��
�2�]���xV�8\ᆘ��%\�;ÿ[��b�[#���Wʎ����.^�|�P���Uh�
V�* )�
F�(๴;��o�C@����*JH�vɉ"4��w.E��J|:�� d˨`u���)�z�jˢ$9#hkS�g��ޯ=�-��M�u�p������CB�lxd^k���H�7�c�*e�aVS+Ѭ�0c?&�4%&�*%Qh�؎�ͭ�ߥ�*3lq�a$�Y%g��iy�4Qd�*DY����Z
sF���'Qp��(j�v��4߭D��<�)��D���N� r�/U������Q��4�22̨ �,��B�������alʠ�U��$�#�mdV�*������L���K&���L��Go`�*G�9]07�-%I��\��Ɋ�F�e�y8���d2�Z�����8�B�,U��
7i�
2
�a�/j
�jB&�����f�-�U����o�*[�C�\qNo}]�Hzl���w\���i	Eє�{�a|g����u�������K2�f��9:Ƴ��Ȳ4��˴U���Ŗ�N��1�Ҍ�1��Y��#�&��S��W� ;%�.����j�I�cP�X�+:����x��b�]K\�A����9��ׄ�c|�l:
eD x(�ɵ�%j��{�x�]Hn�E,1����D�HS�.���F��XZ �f�M��7Tb���Q�]��qs�ئ���U�A�����c�m΄W}�Z����lP�C8��|*��÷�1̦%�7���|��<a��-���k)eXK��C�¼.���N��s�c��+z��4��!�0���AHCn�w͉���V�e�ن��L)p�^�������V[�� �/O������p4p5��h���(�s�l�6��;\Wą�[�Jd�ŝ`�񬋛�F�K�P��i@v��z����HʅV�CO�%8�a�
.�oG����6��l��-̖�>\f;j̰ɸ�l�0s��P�"2����C j�23�iU�|�jZ6�e�b;�=)UV�i�|NRF�3�HZh��)!�@���O�dy�J�vMwQ1�b��y8�.����[魥K A۾0),������b0T�ѐj�)���y�X�eWa�p�.!�m�ʬX����,�:9���i��1��������Hh��4gh��L��!�s����\me,�k��]y���j�%�w��k�����
Q�I#�<-���ByU�^L��.��͓;���3��=�ì��ڼG��pH�.*X�	����Y����T�T����,L`�)Q��MC��7b��2 ��2�b$9sL�<l�(L�)�)�H�6w1�\�#W=�#Df���(��i��n�hr#�-�ɑ4�����X2���Z��> %�ھ��^�h���cj�-�}��oRF�!�2;nҔ����Ls�
p�^����I�i�hB��࿱龬��0&v� KAp����*�7�s��G-�<4^We�3���G5�ě�"���E�!����p�Xg�00�#�26�9sqb�3+�C5fLg ���9�6��(�[I�(N�*E�+����zвT�VW��6��{�=w��Z���D��BJ� ���8��:C��04��`�W�VFj�硊�`�����Z�k��-��@ؽȴBf,e�s��Y@XoT����) ���|(+�ۜ%�6#e˂K����0�qȺ-� �f0�c�T������yOҦw$Q�_9�0FI%�g��^��o\x]�W���b4�A�1E���P������U�X� ����B�M�4޶%h��B��\e���.m|� ��Ѕ��;����%�+��za\>��+�K���L��pP�e�W�m&��ֳ(����e�9����
�Q�[��R�J�H�S��f.nq�$ɳ��mWE�6�^2�xS��A�bP"�X+�ck	�D���"�!���0�D-c]�KQQuR&iM3��Q�\)�֌���"jhQ*�q	R��x�x%�0P��4{@)R����Yf�Ζ k*�8���������D��1��Ԡ"���8bU���
�ׅ�}��Aӂ�n	ٷ� ��Y��Md;��Ve}��iF�d��$�T��d��^�����*�6U�T�Ѷ���;^�%YEr�rB�� �F���\u`�k�	7���6 (%V���1Þٿ�,B�{�*nP\�@h�bNy����!H��)Vh�j�e�P
�V$�����q�-�X{�&VDr+uyY��X+�d���W�0D/W(\�k�o[FS�zq�Dm�01��V{��dD��c*�fBIy(�x��jfu�*J�
�ੂ��
����^M��nR�,M)��.���j6����h�N;4�,@�LC�E��aa�9�����x�6P�ޱ���fv���5�P�G�]|G�t9���F�#��EV�:ON�r�f�⬐z�:����ku^�lB['��3�b����)JUq��/x��l].v;��aL��Φ�6��B�2�a�@��~�Ak)%TK�)��KՅ'm(R�P\l�1�ULBK��)��̥�Y����wip���\�x��#0p�|�s�g�=��Fk�@�@F����a2p�x(�X��$r�0VW*��3����)R��-�my�]q���v��9B0�ͲW;/�&PX��aT%������M�iM�PU#nY���y-z�Jړ��
�)��.׸���bҢ��V#� �j���ajN����[`���z�ժ�7(H5U%�;KQ�Q�X PU/���3	b0E�&�;�Z��\�"¢x;R]:`�\�51!H�lD��ʿ��r.��@]�N��R��;�r�a���5����R'��tμ��7$�"�R��b��P�x�����b�,�cG�.�K<�q��2��3vE T��Ի� RJ�ď{��"��6��L��6���L���`��R^��'D�Qb�R-E����cE���zEL�=ۨ�D)��Z�^�/��R�ҍZ�ɀ%!a,) ���a]�Kl�c`HDIBߚ��zDP˫�w�
JC*U ��7�a�.,�2*`6�"*�TVT����
9�b�r���DR��-BD\N4R$�P�rʨ����V��EZ�&Hڼ��W	`Aҋ� ^o؁��e� 	acW�T"��f���6y�v�p�^�F���!2"1[�i˳>�v��7#|4VT���Ҩ��X�H��+�4"de%k�lp�/P�55�L*�Y��9���bp#�E��X�����W�VX \�o*ň8�U��F��� $8�b�P]�4�Я7�e��k�!I$�H6����u�>,1��<�,T���%���BƔP��B
�6�H��q& ��M*�F5�������}��
\���!@c�Z���J�ʔ3:� ����}6!�/��᷶�5�w$���*@��ɗS��p$A|�~ $E��:9�E�$h��*��D��.
Zս��h�*6`(	 \�1�&�5]+r�"��R��HQz�Jk�S$��-0I+G0�L�
�Q娄�bN��j��(��Q��(!�#c�5 � ˮ�n�&(�(�dxY��1�Y���V$$�RO��4@Ȉ ��s�pI	�J�Su�j��:��.SXdj�ٕ�H��D�.�ܨ"����+��n�H�g�Ͷ9�dSr��"y!Vp@U� w��	۵[nD+r0I U�a�	%$jG!�Œ�`�1!q\s��E/0���h���E��S�� Rb�A���ŻN6RB�Z�!	�ڜ�a���	�����g��Al���;B�PTQ��W�U��V��łH��RH�FU��I��"e%_�;��H �摰bP�φ�MnR6p�*GD%wY�q[�\�?$�2`�.�0DJh��
��b���UEMJ��"� T��^*s@6�\�As�)܀)V©�Y
��E�Ө��V��;QtV�c S.��;����b��dr���P0�.#I��S��H�UTR���(ou��P�+v��������6����7T�,�O��5u$;���Pf�2CpC*�ɾA�����"l
��V��`�%�DX��\@��R��fYMT؋�^�����F��أ,j�������!�����ȫfF!��O/}&�S[(�� �UX�d�ă��R��4��0fH(����d-��P�	&`"�
;�0(Fw:�5]��X��� S�������$GyZ�ndM؍�vF�q6���A�ŝ�J);E]��W)j�8z�m�C%宣%�PS~�d��H��
J"vT]�U�ު2\�4��9a"!�y�f+�FW�=V�
TT��'��B<*s���� ��f)��d��$��)e��5Eّ��Ma8�T�/�ARN+y�Hc��2��!^����c��*����Q��e�,�vn	
"�*����BJ3���f�b((&���z�7�lR�,�B�	(S:���3/�i�C-1,B�K���鸀؈��(�f��e�*��3�v�.�-�\���u�l���+�;�* `@b�飢5=@e�YB�TRJ����	�K�`�4V��]�A4�E6h_0y��Y4��;5`�(3:�P���0��QUv���x>LH��+ٷ����1k�]=��4��������l�(YT�l�X,>�	��̶�M��T �E$)*�1�8�q��H�R�]�7v'3�e��Tt�0��f-&e+�8w͟�S2@$)��q���4$�6ʫ�sff��x�줭S���&0|��a�������}~�%�aK�UDa*!`,*��$ �bmM�5U5o�}�Kˎ��u�u��㫑wr:�۩����$AU�@I�yO9z 7&���XSS`ՀH�EB"�"�B(E ���P����dVD�-J��P��XT�� �B ! �X+�C�}�H���I@*%p('}���7������� ��	� �R@т�*ܩ
   D��R �"� @����6� U�Զ@.b(FIaѴ �Q,$$@$��EI"�HHB�
DD�_��$d$.R�\�)B% D�"�P� H(�H
���}�K�B�$��^�%�T)V,����ll7 ި2�H� T"�V� �I����2>`.^���-o����������~^��0����"QT��3!J�g��@,[�wT�l�ܖbq�'���nl._�?T�8��@�A�����E��H>Ym��}���>Ѭb��V����{9\���d	P� NV}�~��<	�;1#�ӣy�v��[|ֵ��n��) K�ضȔR��- �DcDCm�nG�{_��XOv4{c��,z���u�M�z�L}��6s9	�P���C	A wx- �ڿT\��[��\&�U�d��4b�6��جmĕ��H�$cQd�T6����܅��¾���?���/@�<�Rb�-g�t�]�=���j�[[�����^T(�W�Piꬸ8�e�aARUf�P`y���b&� ����U˚8Cp�qU����Ϸw�k���}5�K�t�s�5�;^�T���_u�{Ț&(�}w]wb�d��ٶ�U�V��ot�\'w�nn��s���D�wEw]�V���}_�'w[�u�1[W]�Y7wR�w:C�r��.���nK�H&Cs��t�*�QD�
$���F��@��j��g�o�}�w�����EX�m���aH�!�_�V���V���'�m����LU|_�3���KŅ�ȩ�%�ҙ	a�$U&Ke@XHWȾĔ�F�TPQ��|$dH��y�1D1B�R�e����¢�{h*�B�(U�$..�HFBT��(��>��T�O�O��_Lo�/��y���v��9���b���=8��E��v|��ubLR�|{i���~�~g߾��O⑄Xy���a�X�����������_F�8ל�81)L���淑�u�u��T2�B�I����йcP��
T�M@�	)-d�R1�l����n�7��_n�`f���)	���4L�����q�䪙b3GC-��.`�/��@�d��hH�Ʌ�K-��0Ѧ�4d,�űsk] �|��lg�E�
�u#u̒F��c�K�=��ϯ�����d���c=A������߆�}�,l���}�:}?��0�n�>ϥ��#H���<C��Id$�;OçO����o?�:<���Ԓ�K_����t�7�XI�F��{�Oq(z,O:Y��EДQ�8E����D���la&"��I*�9.B1� e�� )5@�(ȸ� �D��"`Eㅩ@#�D$j���C$-����L�� ����OY<�>�gYRm�+?BO����x�����#�ߊ5U�3<x�(z#E%���FҖ�������ˡWg�dr��� �U��!s}��$l�4t.�\�뭒�&@@0W�IFJ.QB�JPR�1���^(�$��6�����QD�L
�����?����B��!"AB����\���4D��Y,~ƭfBH�T h�qr�� �(�TT���� @PP��(2(�(� � �����r]l�H�Kd`4\��"傖�$dF@��D2�&�^��Kļ�9jt�����,"�BH�H�I"{����� ����n>6(Ȩ�.U���}���@1B"��!@ㆸ�@���]��}>��΅��zM+�����ݟ���y�.OГ����΄Ñ��(;����=��Xۄ���_iE�.n���d �<��(����XH?*ߕhp`����ࠊ���Bc	&g��G��}{!�q<'w����r�ɐ�'��@xmj@U/��+dQ� R�a?�+�Pz�M�Њ�������MO�w�͢��{ރpt&��f��h�b�� H��|��>l�9�hS���Y2+w�?�3�k�2��D�F#m��l�����(���
��m!�0��u~��r�{��U�@����JG�64|��,�5qdCL� W�|�,���,T�T�	���g;�d<D�>9��(>����)C�G��8}��?e��)�`(�X<�-fG��6$���A^W�1,, ��qn�s?�Ŀ�P8dbe��H2 �	 DF6��Z�����䪿������!~	�B66Q���ȋ�r&����J����X��0���$��Uz0(iF��~�]�_+ey��R`BF����HC"P �S֩@�	x�r����"BB2I$� @\p[*�e$`*�JGP.��$P����2�oAAa?ߨ�1ubY�-��۳������!}UJ�$���0�s�
P�AM� ��(�[ۀ�f�� 1A��+f��H(�?^�:�ݥ��IkRX��8���\FM����JD� DZ�E�=h ��:�p@��%��DCd���2�͋��S�AR���:�&����2�-��1��H2H�/�Rƒ�
�6�SMڀ�`�CO��5RBN�B�C��$�XH�2I��@�FqUC�b��mT�n�� ���[���w�"L��xg ]�٣��M�dD  b}� �h�����%"�\
� @8��Py�o�ܪ�� 5B jc~$"���ۄшc6�cd ���*a�YPpHn�v*�ttT p��Uȅ��� 8���o�2N&*�"��,vh���o^�2�`ͻ�u�8Q�V�z�c�F�R ���\F�5�
xlt[� �q1M%�Uo8�8�@l@؂���� �Q���BD�OP��QI	�+pa޲) ��^<$�T����p��T��b��, X	�!�cˑ�g��+�	��6,��������ݷ}�mu� ���t7!�nn�&�֠��s�t����H�d��9M���ݶ��&`�,��8!��G}�r�ψ�B�3�1Q�\@2;p
J4�F?��Wj�z^d*��DC� �DBp�� �@��Q2@�\M?�E�����6f&G�2 � �*�H�#��|�5�oǆ ��C
u��MM�؍���m�a��{��<��:d�0'p��˗q���H�D1�mu�P G�م��c�������{��:A7�`��Q � iX�7P+���Q���A��g��ڀ ��g�!T6��BB�����A�[�D	ZQ�2�/
	` ��~@)�AN:.
A܁�����	1ZTSXV�%XK����
[�$� ����\� i���� � m���Z
�ze��m�4�}%" ��n��i��h��V�H;nS(���a]s���O�D���N.��B$$X�.]"�ny��/C���x�@�ρ���yzm����Ht���<9�v�D�*P�Z&�B�DF� �qAjƘ��Wr�*��(�-�) 
�6� "��һ%+8a}�8X��j<I���9JI�n�Q@4f �	 E H��k#��< ��*�a,�� �S�:z��S��|� Q�D�!�̡� �,���,U��K
����Z�r�!�B��>�(
7����Z)�!F��YL�@)�]�[^���
5� @ᰁ�@ b��f�(9P7�|�D���-�Ex��}P�ou� 5��_���! ��(���j4��v�1���_���X5�9�ܠ�?"bVtq�j���#!��]H�E8�"����4��'�l��@�����(
z>��[��%�)!�6`�ڛ�suQ$��Om!�`�i�~�mx�#ǁ�}��D8�8��������!g��_�4{Si��>Ϙ���U�@�'p����_�OC�G�|�1r�{ �r�T^�0�\�%��G�>-]r	�v�Ժ���]7P�_@g,r�1՞����t�v=����>��=%"��}a&��Їε&˗
�D5��H��PGڑ��$���. ��H{���Y�,@I����7��4b"E����ѧыq�܅���px�x�D6�I-����D�������Jn͏}>��|�§O����q�?'����,�D�N������������+>g=m����m�����+���÷��d����M\�9��ڽ������L3w��ݷ��m�A����x�ٟ��/Q�'m���~�?�x�� j��O���I�����������$������{������J�y�ty�?���2����'s�?����4�6�O�a�w�Z�&���?��K�x��,��'�!צ���j!�'&���?���ƍ�߉���1������+m�׌�q�\���/�������۟����d��Ȗ?�g�iy4W���|K<�|��$<����}��&�<���_�_5�>h:�r���]W�W�^�_�k��b���~/�.�<�M�H)���?w�G�d�F���'l��_�I��X��>�o�C�|<s���Œ;�>4l�H3�-����k�4����+.6��~Ū�7M� ����7��3�����-�������Ơʾ�/����\��%msV:��w���p�n����������'�?j�����o�?�?���b{����������g�����~/Q��?i����q9���������?���!�8�DO�;��ҽ_̇R7[��$<��|��s�Ok����?/���?�����>���������~O�~�f�����j/��������������������}/�����l8�V�O�o�������}�*p��W�w��X�w�&�W����p}?���޾�?��w�E�����m/?������l�"_Ȣ/��?���E������'�PoQ��������{���f���D�F�����ɵ����>[��*�������4������������.}؛}�?*�?G�E��>S�|~>�1~</�u?�� 3-���Z��g������}��k�����y4?_�����O��Jɘ�J�k�����]����s}_������6��C����~_ڼ����QȂ�����n��x{@<p_�K�_��%/��=�s�VE@��5Rw bH�5B��r\P8@�����ަU�p�AK0P��vd�@_|�~ ��S� s_d$%�d񞪃ÄPQ�r���Ԡ�C(�|x'j٤u��B
���'�<�������������o�,
ZԆ���z]d.O���eo^O�}x�A��xe�~� ���z����҈/.uE!��2�hO��^BW���!��G��$}�y�@A�?����[���ײ�:���/:q�:����Gc�o�O�޸�~?7����'�͛�ї�iid�>~lݍa��7�͗OT�:E���-�Sk���D�p�YJ����؋����Ty��rA	$�!�83��w�^���\bv�ᄔ��I�@Y�.�](��$�]q<���E�/g�?��<I�J9^�q���<to'���=l��N�KBAP	�����o�gE$�H3◇hCH�)3� \6u/��x��!$��`��}p�J
~h�
�vA	�������]�a!% �����f��b�O�Ѧ��p��>���fR)@D��җL���T�������A࿄(��T�O�Wu�q��V'%�T6A`RE�E��$D �PB�P��D��,�h��� DF�q�4W��G���\� J<7mϥ�{�U [���7#r�XT� H) H� Q۞�l �.( �HEB>���[�"-" ��"� *EX�@�AH�@X��� J���(o�UVX�_yb�@,�U�EJ"�T"H�H�H!H)`�T �t�HE�d�4�z����kj�O��nq�'\���.]9�)�9.�׭�ߑ�Q���O����?A��鹻��}O���@{*]gk�X3����}���[����&-�O��~���z�|��_!u�%����.��GDx�
>A�+��	��B�?��jn?���W_�Gs��A��SQE�d֭�r�s��a;$�\(�@��[B��׀���Yh(z�LZمb���0�!���
�J.g�t�t
]!�9Hֆ/FxEAs�2j�Z"P"H $ AXAX @@�EX(D �P�$A�@
" @AXR��cHf��ڿ��Ѭ�K`��kX6��hQ�	�f���$�z�Z����7�H���X�s�M��Q|���t����aX��6�a��>��|-�:�R��6�8��>L�:��2��^P�^8�d�|Fvl-��|@�½1R)'�J�5Ys�
��7�"�-
&��b3�ߋj��U�^��(8���5_?
F+�e��5�/+��i,���Vb���t4�mƴ�a�"Ы�T�"@&�o�o�����M���ML��� �N�̱L�1��Mއ7YÍ���.'+6�v����HK�/,���q��zM^N.�ĸ[R��!\oYV9���{K�x�6�ܽ)��FJ�J�Hl66��,mv�Ƹ���8|��j4��.t�� ]`�dL�\�h�X��������5;Ꙥ� 6y���O�-�#8�xR<Z3�q
2���~���O[o�-Z����c�Om�7ԕ��7#��u����,�;��fj�3�4�mZ�X_���f��̶j3�k��m[W���x���;K�jژ�xz�L�"O�j���=������:�R��o��������[7j�h��'�_�q�])�WU�v"�����\dXC�]w��G�q��^c;�}N-+�߈�(s�{gs��8~܊��!���te��y듎;kp�ߘF��o�=f�[�lY^��m�jw���|ӎ���������h�_s��CK�Ɠ�+}���Q�nNZu!���n3-�Ϩ���;m,�y��pU��%��3�1V9�w��re����/jʝ�N��zv����u9�٥p���i,̙_}��xq��������#��Ya���4������ߊέ�ݚD)��)��8�������n���!������m�e�{��g�ѻk�����o�8��v�����^/jq��mV��+�[lil-�},��2��*�#V(( � � �?�O�x���^|�O��������ō#��i��?>�e�I7W��������u8��]���V2�v��5�;[׿�CKL�Z=�!�|��^�ټ�����}�w��kC�N#*F���C�mh�^r:���=�xN�}�38� ������ϭ�voi�ݙy�3J7��Kv�S�m�u
�ǯa���b���g��q��z1�zw��Ĭw��q�n���5�!�uX����<z�:����Ubuߥ�1=����V��;󎫏T��]�OȲ��|Z҆��5�1������AU�߹��Ng��;k��Yx�G;�N���o,���u�M����t�=�.�׍���Q����냽kj}[���<vϷ�\���w:������i���ɷ[7��oA�c�g�ݟǋ0�;���7�KOm�����l������6�}�������=��(�s)���<w���6�����˻��W�-����p���a��>)���Q ?��8�`\EN���X�,#T�"��!%� D��@��D��������@��� @{v�x�[����v���6��$}~���~�m�����>�o?oM�7�C]Z�W��������lv����=�&�-�,���ϟ���[�{{g����,={�>/���>��ϯT����?;p}��{v�;����A~�/E�zW�V�zjy�����>e��ǉ�w�j��o�����Ag������[Z�~c����OOߎ��?o�������m^�8�k/��Ʈ#�ۿ���y?o���c���=��_#�~ͥ��3�r�!6�0�HyD�$qQM�!'p� db�(���G�/�w��٤Fx��y�|�����q�����ۿ�ϴ�ۇ��3w�C�����^[y���_��<��>l!��:��Uk��
����:�S�R�k��K��K���L��K���o��>3���8�f�^�X����U��W�y��|϶������(a=��蹨�;}>|za�q��v�?�m����}z���{�Ǟ�:Y�����F1��t���7l��}c=���{ʷ;o��;��>>����K�s)y���|�^�����ckߥ�oS��xo�������Z�[�=y��;[�:�n�J�k�Ľ4�\���g�ݾ2�h��m�{���'��n�����d @�
"E(�_�=�}���D|v��%Z���R)C������F��P��aQ�8�۴[��������Y�*�wz����7Ϗo1�\��ُ��.ΰ�TF���������;����걔�kN) ��i����Ld�}�Uv$4��s�8C�2YG'�M��F��Rt��H"d��~�U�aeyi��H,e5��s�������9��K�`�m�y�f�����H�зi��T!xSr%MA��E(DU�RHIuXZ
�:����	�����ow˘b6�#��<E���v�������_L���m��K��y�+�dg�g������
{1j���7���~�����u�4����v�c����m��^�C��~˟��2j,���iÛg��O�H�!S%�L1Ʃ��!������66�ЄF7��;�%�O>��g>� ���6��l.ˊ<���D�����yf,��1�މSqp�TED^%�`��X���P\�_,�X�<�H^E�H�8ǕNU��b�%��fH�|�����I�����ip��#�!c�"@s�)���d0P���P��x`4D��ɤ�6�5�P�t}��#��6���Xu��?Zp8��{�����Lxb���f1 �%�|B��sc�E�Y8ux���HJtbP��iGKQ��(TR	�>�Γ��$�X��>9���c^/�/� DD �O���Wۿ�5��n�A�����M���E�y�(tW,�I(�-�k�' PȢ�ԅ
��*�2���U����u(�[���z�[�����ǟn2�=k����,ZFA YA[|�J�.*n:�l�����3�r�� ͼAs�*$4�P��u����S.�FHz4(BEV�O(��¤�ژI&X`����2.a�Nr���`M�~`[KP�F�@�|�Q<J� )��L�MX�����$V�Y�2yȪJO1B��#fХL*�2p	jE�@��������P�$�*��BI1�sl˓2�(�Ӧ��΃�/$�
�,@yRQ��x�Jx�%u����)(� ��i�F	*�0�L\�sKbu�("4��ЛTCA������an"��Nj�B\ӹ-0Z�+(�|���)ä	C�q�Y�q�M%� 	X��+���s�F�R�4iB���؇��$��)���/"�#;<,Ѫ>�k6Ӭ�$8�/��!DU<�©���PH�#x]#UW@Td���`Ԗ��֒d��b@3kF�$.���`墰f5��YHU� ��(#U1�9!�5ɀ���0���,��X�;Lzn1�Y���c=�
�[���e�q�G*�CK�X���s��.u�(���b!��LG���������u����v����x�~��~<��A���U0�BM�;hXǻ"F�(�1

�*�@uN���D@�Ҳ����:�ҫ:�ۣ�)p���<����L��9q P"���~Ku�?O|�����s��͏����-H֝�f�P���p������U�:�:c��g� Te#��1:��j�O�z�o��w��?��Q��>.��H��o��o��Ŀ4�"�3VK���������p�ꢳ�$�,2K��Ȯ\��Ld3�1t�N���Xc>���@�u@N�9D\�U*T�!$�sMV!Zv����,P�I��M��^A�!���K!��5TJ�����u2�T��r����NN�W�D�`�pH1�`&q�$�x�Bs�I2�X���>��"Ziz�_���J�b��L�PJ-��$�b�E�(�O8�EG5)@��' u��d\2�1d�S�M��5W��"f�T��}dOJ"6WdU�Y��!�E���c��DH�L�̭ʠ�A4����Nǅ%O`�g�zi��h.�".!Jjt�%ay"P
�b�1��$k�6*ІY��1�hc���1@�8���<5�
U2�,ԽL�8+Ⱊ�
r�٪*y`�X�c�>��D�9�Q���"�"�ZG-CI�#$5<Ȑ;�Q	S]b�ak�k�>B�H�d(�5ּ3q\,��!y ��q�$��d=4�I�M��68%��He��'E�֥4TJ��K�=�8+* c� (Wߙ;�R!��dg6		�a*(K� %0��QJ�Պ3%�v�	�ʠP�T.a����ˮ��G)R�NN�T������7�}�E�2V9���5�Z<POQ��R�Bb>��d��1��4�"!s
���L��4j�ZU#+p,��8��I��+P�����%�R�H�Ի�=�=J��S'm3�B�J@�Q, J9���D�zY)ɸ��8�*���j��y��l�P�A"D"@ �T Q )#�H��  �-�)�@�������*j�,��ӿ�(��jK��
&�O�x��u�IT.(��2f\��눤����ysR ��"��_H�����V�	K�I%�!�P�^���-�H�A�aK�l��笡�T�`b5B��PH��A��Ak�IF,�e���T�'�v.����Er3<"Q�7
�N���U$���uj���v(�y5�u��j�072�V�V�%�^T�]�bA�]|���+Ub+0�ΖB� �f��QI���v����Q(��@p�!|�^��y�Zz���D'��ＳN��1���6�Ҟ�Z
Oa/TRc�C��Y/,� �v�4fc�4)^y
�* A>`�a��0���ځ��R�d�O��ӵ�(R9t�kQ�l���$¶����vS6���`&��N�G���d�p:2�>��(�(�b�>�9��-�PODfPL��y��zy��@����؃3=T�m�Nb�J�˧s��6�+�h�F�E��B[.�Q�`uϑ�C	���܅�U!נ;	��_S�LK>�s^�w�E2�X���
���d��HX��)RHFx��B#m����	��
����j�#;ޑE�A���v
]'q�X��6��"���~��Z��EVN&�B�� ��Y^����b �e�R�t�)2dB�p�H��<���A�kUr��Y��lR~�H�9�0z�x!EB��=�֠��IS�[����1��f ����LB�M#�tW� h�%S����X���U�6�]%Ġ9���(m��2sl��~i�u �sI���B2��P"p�JIU��(	a�L%�Qn�R�B�UAg�<X��V)��%EE:KTh�P�R�Z}S�53��jϾx+�f�q��¨���v dv�����J5S�g)���a�K/��/�۟�����ݛ�F��x*"�� ��v�գ3D�S5gх�XHTn�K����d`z���^��-�(*8U&�ȷ4'��6i��	�7�hM�P�TiN��^�a�d���I"�	TR�vt9ݙ����DV�^O��Z�Ŵ��� �]E�2���E�lՠv�*b���0��Xp�,����`~�K�<0�$k��
Zq@ZW�,3��.x1T�
4B��E�T��Ul��%H�
��0�ħBLY)��*��{ ��ѷ$�L�-��o~��L�D�ɪaj0�}r(�(�(tf!�26q_;��\Ej�L�0�"m#B-0�� ��TcF��a.$^JK9X���A�Nd�U��	t��x���L��/�D�T#Um�*����'7��&
rS�@@F�%΂qŘ�^D89	�8��ヴ�M^�+L�̡ V��Q��y���R��3Ӯ��S��*���Q��`e�"0a��/X��\��*J��Q�f,�s0'6�Eڍ��+�K]d�c.g��|�o�H���"�QXu6--�(�zh��莖�p)s��AV���t]7n��ZE�$G�* `U�钐pp<G̀Ī$��]��*�4&6�1n9V��LS�JUY�te��-�X䫚��F� �E{
���4��0r0Z�ӎ��\Uà�e�*2Y��#(�R��j�� REP�Le�&��hB߀��D�Ӯ�S�M)�M�dQfkp�W&��M���gc��U�H��X��6K^	ơ�Xھ4Yj�J�Y^��_GW��(��y'�zy�iM4��h�Y��:�4|��ٲ��bed4�U ɩ�����J��3 �y	P��;���m*�bxf)r�v�R��)����3��$jA�Xv0^%
T
`�Rh��k&�22*j��+D}�Bܱ*��/m(+P�.S��[�=����P*�tM-E+")�<R�J�U�0��*���A�Ȓ����	�6se��u��[V&��Lx"�ĐuO-�Q�����)s�՘0Ih|����Tᔒ����v�
P3H����� ��cT�� ����������H�)he<�f����p�G�اo���5i.�T�z�g8.�ǜyO\e<}��U�2IȻb���;����,� tqRF����CM�%�*��{�-�ұUI=��P��E[�rD0��<B�+�<B�5n�D·r�;�& Ya��f�F(({E�.�Ɯo����+��V�3[y!((�Gq���I��VB�G+��Y�Ɯ�ח���+:�}r���]WY�`S�\A�qnDY�X$�"��٤�E}4���^��~�Y�ѰxiDU0��˥�H�T�#ܢ0d	��k]r��}g���j�k�%���i�~��"H\�3B�ʕN�RY�ۜĺ���'�-�m^�8N����|����DrL�3u�>V���S%���iBO0��.�fy	V��Q[xk��cd��D6��Ր�.5M!Iר1�չ1j�L�*�����GlG��=�#Xx�V2��4p��E��+��*,Ђ�����d��!x����T�Uh4$=�
�B�A�S{p�U5�[��isaU�.{�?�[c��*�!�Ը2���V�(U�E�=���D�J�Ez�2�k����U5�E27�pf1��ؗt�ь�����ֹ{&�*�FL�Lmk�k���L��a��.bst�jSIN�ʌ��Fj��Į��l`�V �H� �殚|=Ec*��労YiqJl
2CC�fz�Ƣ4�t\W����4��EL?Z�e'��� r4�e�[UQ,��qe[�T()�ir�vJ��KQd>u�>�AՅ��'&w�6�5�*q0{�j}<S��!�,ƈSW��\��-RL`�#�]p�a|������}8!�gQG��E�Q5��QB"���8
�
�&+-+veO]�T�-e���aZ@�FLX[�V�J��G(wJM�E��3"�#'j(�%^r�]-�4�1�z��lR�9�Rx�r����2k��l�B��(�
�=�Z�mc�=ݸ�q�F7���������x.������!�T��MۋjRǄ��|i��`�P�α�[<2h
k��BV�O�%
m�a�ru���i�w�8n6p�>�6NHWv�޵@<t`{r5]�@�g��+b�+@��.�6V��	樉� ����h�e(���ֵ[��N�s]�m���gZ�W,�$E�B-��1����Z
)1�[\�sF��wu�:�3����
�c蒋I%�*:����I�DV6�(�F��l�n�V6��\�rث�.�F����wv5%�Qk]EP� ��#",�
C�{���?��^����ϧ�=�a�>G��]�FHI H0�I$$c�D��"AF��j+h�֊ص���6���mQ��5F����-l�6�0-�%2BD�fVV��6�	(�MF�LQF�56 DhJ֬V��	$dEYP!5�6B6�kcmLd�!DYY$IEDBAQ�$TY@�I�$AP$DY$I�D$ �E��FDY D�$Q � DV@EA$$RAdAU�F@E�VDEY@ d@BEBE$A(ڪ���kQm���@�UP�IBD!��$Sf�Ͱ" ���
,%¯����������{����y�������7���y���?��~��<�_�����ki�}?�����7�ӹ����ug�㻣ɀAa@����334���"a&��5fB34�2`�ҁI a$�B1� i&���,�Z)��1$F��S@�� "dL�%�����A��&d,T���V �,ba!��Ff ���$X�Aa4̔�E��e�Je�12*�($E�Q13`ș�! ��20H1��HD�I�1@�@�d	J@X3&k&E(PI4�HB��&�#4٤�	M"Lfc,�L�B�$�lJ�$A�FBIQ%`T��	�$�����E,�`2~�o��|�?�z����\מ�P�@"��w��w����.3�~�������=����m~7��_k����r
�e߼�a��6y^�����%��U������>��/�~W��M7��y��Q?��/��o��r����u��g�����{g�� �8S'����{�~���ū��U��w&��V�Xȍ��2���B?��jKz�'L`X)��M�]�-�¡�	D�:&*xY�� ��d���4��YN������I�>��6X�Η�-�䞹D6�
�D\��������� �[p�-�\�U]��9ZZ"veS`��̎H�9,�m��\�8�����sD����'Cb+��G�1�r�A�#��,��,u�@���{Z1(�TES��Sz�R�zg��ή�b�s�Pua�&Ff���6��H�(K�������
͵����3���h��[-�U
`E*RIn*��U-�2�+�à@!3!@�lQ ���T��u���ЃA�${[.�����LgE��@�<�t�<C��B'K�.n��}�=��P������A��BE<�N�n*���qYfT\�E���Gр[
�%����7"���U�<4��)p"{��t���<G����z\��He�BǊ�bu�Q�O����
�2^D��̊\���:�I���Μ��<���t�5M*e��y%^2=y�@���a+�)fi� �[���܅9)ё�G2Q��W�qD���s�Heb�Kӣe؛�ޝ�4��ܒ�����^*�f�Е�9�7(;Z$����Dl��e��X�\��Lu��JU��:dv��L�(� ��Qu��i� T�s�N��\�t��k1��a�o=��R���>����W���PXX!)%���[�b^&�+��`HՉ(7��䴥мG�q�J,l���7I\d�"�{,Ԡ���Yʗ���:*^���:�f�6Nh��h5�9�AЂ^��d��o�U]���K��I$n#�$�X4�J
4�������i�(RA*�������@l�� cm�[m̕�|�1Y�J��zVN�ҥe/e`���2dU^s�d���8����"�U\Ԡqo\xy摰q�����vm��#Y����u6e;�Πe�HS��=��=ӧ"��_��pS�r�M��[�B�!���@��{L]�۶���sK��L�j�4o�!a��z�L�ܴ��[n*�d����z��C<�3�?X�&i���[�Kq!�L�l��|`�U�g+�����^z�[��Z>��6M���<_t���/�r��J��+�߳���AM�Ia�󭈿�(��+"�RI�hj �<��t�>�=�JE�$�Ȉe�[e��mj �&X�W���rL���9eA�6��r���cH�背�_�
I���rDB�&{�@�IB�"
~X ��DIAU�F@UdQр �"��X���DTdT�@T�E* �")"�"*�� "�#h�%AS4U4�H�h�DL�$ACȀ�Z�I4"�TC$	h��*#� �0��AKEo����$T�FкRBE4�s�����$`H����b��L��0�����������������������������������Å>�=Y�0r�m�ҭ`@Q�{A  ڂ��<   P �                   ���                      AԐ   �    z p
  I
���FU0              �D0	:`[����b�     ��t n =	 �p   � � 
���(�D�ءB�
�(j��      ���Stu�'     ��$�5     �"�ɀ    �%$���  /      �*���   '�    � r     p #�                                                       �  ^     �0     �z�:1��a��&� l�D���H%
�H�$RT��
�(J͠n�v�kZ-t�T �)@V�J(��P%H(�%T ��
�	UH$���T��h����P�-ǐ @ " y�����a�H������0` =�S@    ��   �%  �L��)/�๾��@	 �� � >�(�@�(�]��A  P@  ��$7,
 F�     �d[{��U?      %0!<�4h��a�i���)�O*o#)�	�i�Jz=M=SD�LM(&	�F���5dz�i�0=Pjz  @&B�J{TzM���ꞍOD��?T~����dђ�~���@ h�5?P� �    �?
H�S�   � �        @        4   �H�"
��z4�(        �                  $�J(���4 i����2 ��  �4h 4�h    h   �    I! M�@�	�&�@�d'�C4�4 4hM� ��`i1��Sa4�d���с�`Q���|� ȫ�(C����V[T�������Ě����<��9��Гf�u��'g2�����ۚBq�C؞#�����le텮����B��t���o�n�{ޒ�r����z3LC�<G�Fq��є�i 3��8L��^����-Q"$[@n�L�P�����������z9�s����a6�E�aC`�&)�~]6-�ʶ&�@�0�����UZ�h뀉�  ^l�Brg-�8��{u�^�q�痛\M�J�UV���~b��W�_۴(�Tc}_m}�f}�}ܤ������2�?(������	6�������㭛���9z�E��x���%�a�f�K�|�A��l<,�q�L�R� aaQY4V�K�}DCl���'
x�>?k��<��@6����Á�g�캰������_V�Z��ax���
��$Q묪 x���uRB��<EW�;��nt4c?�Ϟ/�����a�|�˚�-��E@�(�۸�PTKc����O�� �I$ %�TQ�H���E ��:�Q�X�$��!>��~�}x�~�~}��M�xަh^۪3�4�i���1:ƙ�)�fI�4D ��bg��.�W3:f����,<~%����J��He)�^0��IĖfBR+���}�i�t���l`�$�"g�Q !G=�}#i�L�4��30���i����B���M��U(�RM/��6%%���9���*�а}S��C����;��ǲ��fg�cX��\�]QD"m{f٥	9�����7?�y��iެR���Y����RR��j�>�G$^�{�q�0�l?�1��,#��,!75��u'<�\b\�Ĭ�X��{�_1�^����?D$B(�T!(����30?�o��bV�@���4WbC@��f��׎�9ZχČ@���܁�`�C�M�`��:Z��M�bs�4�˨jh�ǅ��[���VI���v�#���M�%H-��`.Ypj��x��H��b�[�\N��at1`╾,�X��<�-z�P��P%j����[���a������%K*��g�M�q0X1��5�0�0��l��+�C��fB0�|�#X�)30�� ���`r�	`b1�b �0Ej��;�iye���VΦ2�H�	��o���D��P�C�0 W��'W���~�3������ĉ��ol@��٢K-{�F��{�e�'�s��dJ�%�˨p��~b7�~��_�c?�jF����j�ߟH-^�W��=e��(����F��r�}���5����j�b�?y�U����������������VS����������b��6"=[	�����x:�c�����?�EgE�@��/σٛ^��A�_�������WW������#�f���P/H{_b7zn�ݢ}�ٖ�nT���W���{�K��~������N*,߹ߕ���E%�����Ҏ�~�J	2����dǳ1���/��o�
��
���"�r�5���aIE�-Z�r*J�?���Y{��U�o5]�o�M#�n$���];�R�#��<�׳ф~�2�I§��U�
B��G�l����P��~0�v 7` n ߉j�C1��.��hl��  �DaB�� �@s�6 Q����_�[Bl1e��b����5�ؐ~t�l�H�OS���0S[\��h�1 ������]ga���hMKo����~p	��Y/ƅ���*ea�U�D��u�vns $�m��H�H�	B�L5���{۞��-oɱ��H\�5Q���i�����[���W3�<������G�r�Hz�!=�]
�? ݭv��ބ�J�����ˏ�);���We_� @N������8/֯l���_sW�q[�}N����jߠ��>���tw\�k�q��w��sI#;���K�v�I��f1Ŋ"�FH:�-q���MWM��YSW�j�yk���k�� ��y���kn��Ꙗj�֤�ous�<�x�J�흥�]��]�\�܁YH�c)JPec	(�6I�&f1�B��$EQ"ER ���b�b`F�F�)%�W�������Km���A�%�BR
c-���$*E�1$��"�b� $��T�#*�)W)SkS(U1��L+2�qiKm�`�!��`��*�����7#�JJ`D�q�V�B"�X`D�bd`�nX$�j��V�$JSF�VJ��F��Z4�$(��LX�	V�)�T�c-b�1�24����d+�VJ%)a������� =���B����t�P���1��U��Uȩ,�ڙ�mL�!�kB�m�LjŨ�J)��i��d��:Tl��EF�����I�j�E�&c��V6+IQ���߁�����6�+ZTʈ�O)�=����� .8 �U���w)�uXx���&~$"�T`!V(`�:�*D@��P`,P EF �F �R"D����vv/m��m�>Oa�� YNx"y,X�q_� ��R���{���P���Q�0 !D	�K5��Z��ʩ��@E��nu��% 
���nEo��-�;�p����y���L��W��u~�R��(�I�w�����_���O�5����%�����o�ƛ�����s����l/ܯ����������~g���������e�eG��������S������磊��_�p����#�.n�_�i~g����0}v�//���?U����?���TA�����O�	��������͎]~7�gM�����d���7����k�~��/�!���������y�������������������������u�^!�����|�~}?Г�������gǛ��_��:��+��������o��m��'�.�]���5����{��˜���xm�\Ѫ rb�0T �����.v�b�����u߻wm������wM������H?��/��}k�ϊ��|C7�A���;_�S���'��]S������E�|'��g�����-��?�=W%{ϭ�����$��p��H��}����?�����EV��X��Y��7���b/�|_���~/�G��ϋ�~�~U�����������+O��?����~�+O���`
#�[W���G���,c~��e������o��ry[�k���8�����u��k�<;��.P�x����k5~f�QM�V<Q����R��
)�"d�;�ɉA�b�"��|�â�&��.'m��~�=�l��l��Ke�t2���Mh]��[N��TP�S���d��0����`@)~��c��?�|�Gv��@�`c����;���0���r��JN>+>�mb���ݿ �1��^z�u����@�r��>}���6��� 1���zϛ�r� ��B3;z%y;����.���1b�S�7�@�1�`{s���.ɜ�s���. 0 g��׎l�\_�@}9i@0c  1���q8N>�_���4��`c�E����u��^������[k���&����N9�{01���}L�LW��=�<��|����i8Ιvw�H���`c�K>O�M�Ϧ]�&'.���/Ʊ�ǖ���z7�u:��o�[��t�/��Ł� 1�[�����M:�Wk�ۆrk�坒�=*� �yro.~�cί��6�����7�a� gN��]�x˞tG��Zb cݯ����.]���#����"�3��  �.:��[�w��� �C�ݻ�g�],g���}���Zf���1�q�̇A�f�L?�4>�<z�3�<h�W:�tM+�;�!�c c�u�2V�]m?�~�쳭N\7  `c��으�V��*�vݎ�m�8TD��_��)�xŌsYQ��e����?hoδ�U�7��_o�������Ct������=��L�f��0Oצ���pi`��kRLb w3��Ǫr�f`0:��Ӧ��d���O����H<�����N>!�Z�fv` 2�ʼys��sj�~�%�b�8�>^��Y��� `c7�}tߥ14���Ř� Ύ��{��������9�$l0
�'z��c;B�u��ڷ�q���ۺ�0]�������"[��{�ݵӅ*��DɌ`�La�޵��� ��g�喿f|��f�ǃ ����W.�  q�\3���A�C�+G���l8��001��O�J�ӎ�qï����~E}���d��S`�T�hl&�c��4q�p��T�o�
��`0�=;�G�ό��'����noW�޽e������ĝ�#���ȶ|u����W�	˭���1�ڑ~-����ϻ1���E�~_o{���[���w�Q
}m��;�:�=��%�p  1�o]��,�����x�e�JFN�Ɍ` 3!�)�����߃A�#�>|���"�~H>5c*�����FY�����݃6�c�^_�-��Ư�]��8�"<������lw٤!�Y2�8�<��;�y�ָݛ3o~�k�c cr�.�niƱp�gr���z�h�λ�j�����ǰ�o��;GKk����v7Q��c2[HQX0�[���;�?.��p竳}_�'�U��&0 ���w,���E�W}�Ӭx�@c9�\xs���Q��l�]�|>~c� c g�//oҏ����V�An��3±��c�yٌ`c-�<�a�֜4����ͮ�:��.��ƾ�3������G��` �?�c��f�i9-�ꔬ�o��|��|WO��Z���}{}9�01����kY1KY����ü�(�zq���m�� ��>���sU����>�M�{�o�)�����@���􅳦��7v��XڽRm�-����e('����|H01�H�;ח,{j5�%��]�0 ͟���Z1�v��S�t5����0j�J_����Y�s[C���13�d#�y�������ǖe/v1�c8=��9D+��?��ټ��c��f��T�p���k�Ja]X�1�������-�����:�J9>[j��+zzO���`+��^~�߮�Jx}4^y���q���  �z�JwÚe~�]�ڲl{��M��``�vf�u���K���1�ei\���M�gѴ�(�zȅRB6�5wm.��ț�ZJ��2_s�'��5J���[���i:�7\��E�Le!"bij�%�Bi��>ͦ�D��h>3��c ��9Hd5�%,�Js&��a	Kc(_F�	�t�l.���sK���v2��Vi�Y�����Y���v�u�a�u�K��ő�V	(&6  XV��k���b@��˽2go��`�f�8��l�	I�N��z�-a��*F&D�4HX=�]�$�^f���el�B��{t�����lI�8޹g�� �T�&�]�c�獝�Y����[��c@e�;R�N�B�bf�a�Jm�j-U���H($!��6��Sq3e��v��N	��hR S��,���6��]ix&�XE�NX��AK�twZ;{ip�H�L�J8&�&��gj�ܵE��نV�S�Rz)�f�;M���Moh���nM{`:��l�W��rZ<��Ƙ�" ���Ѧ�ú�˽w��2��"�R
a7q	��։�8����ԛl�������'[X��1CZ�XJD�R±
!�D�y�sԶX�!mL�:��q"bC�� Psm��KA&��Z$d^�;�t��iRY��QiVi����Ҝ���i4�����8N����Iu��k�40�!Y�P0g�B�^r�L�����j�4L#�0�pݡ�e�r�b6��H]�:�݈+Ų0��ٶ]�����a^7]vĒ��!*�3l	�5�#(��q0"NQ�R����m���v7����w����0!"�֚�M�VZ[��w�)59��@�����!)���o.��p�rq��r1x�e�(&�%!
DͶb�5r��"	��"	h��X����@�e���AŃ�%&��f�@$�FPҚg^��RRٵ�N��_u�W׉,q�1G���[)ۡq��)5`@WI��6�M
����Ze%T`�])49t�]9�A�]r��&�BX))z���,���V4��63Mլk���3�U6�N�ٽ��eMl��������ZĶ3�3�����	2Y�S%6�EB��K�Mc(������4�����@$
�z݌vl����v�����#	���ʁ�YՁL��C5BͶV�bdJe2�'[CM���X��S�� ��H�i�-�-���k*��G6� C��2���;��,r��F&�7�Y��B@�qf�m�˵).�e8Ƽ0 �.�$�u峷w!��'Veh��6�ì��dp�3u@6��w�%8���4��c���(��M,0+o�L�Ӻ!-�XX�����ve��2$�㥽�!qݛz��]v��cN�ݝ��'\h��ԄD�9a��&����n�ᨢ� 8F�=�S��]Ƿ��Ύ��T�%
�*Kf���'r�#D.8.�u��� B��f��WĲ�S)1`%�X�_׺��8�t@2S)y��!z��r�͔z�܄wf��wM.��*�L�� �!ٲ�(b�Jm���:d�\Ѩ@��p&�v�w��2�r��	M4���L��N�Z�1�^ڶ]`/��X��,�r\w[�<g����r��t�rQ��R �v�J@ۥ��^��HA" & ��r�Q��Q&���Gw�5U�ð�(r�H"�ERi�!JR� �m�h�v�;��"m�)	u���L�=^���[�d|R�$+4��D��:Wm��l�hN�<Yx��Ȕ��IDz���UQ�@�J�B��*&�c��Gu��ͦ��SsV[	������`i�a��Wכ�G[��]�����o<PT�aeҍ�]2�t.����!�����N�vu��dKڣc�*=FF�FV�3KM�m�&�Ix�[x�B���t��K�u���FEX	ŬA���`O+�[��]��
γ�ʦ��+f���"�uh���4�Iz�z���'����퍌�D�@mb��	��dԻa�����CW+����mOF���$�|g�Օ	|�%�fc0���)=!��,j}��;&B�5�m�����ɓ$n�@V_YriT �{d��z�w&L��$	32L�vz�|K4٥���n��� ��㄁�;�^3��H�S��ғ��"n���"X�UX�R J��d"^wYLJb��R�;w*tWL�D��|M����%���aA���fĚM�c�k.x�A�m�]Xv��U�l����8��4ꝭ�q%ؽ:2��W��'`�ki�[��`p�6��u٤j�gؗp"Dά�Y`@��v[B).u���@&��u-�Rp�Iz�_�<E��-��%���Y��HJ:�,{���"HA4�<c�_m	\a &��Rn�p1`I C֔#�H�\t��J]w�����8����iHW6p�ť�+�l#�(@��޶,vMc/��4#�d!��M���* g[9ۆF�o0'Bhޛ�H�:�ƒ��Z+�u�c;�X��R���e�Mp W��w8�s�ID�N#�f��Z�	��J"*.�) �@L�m��ܔʻ� Iu�g�Vؒ��X�H��3���4�S��އP8�.:��vȀ�i�h�` ���{g�v���f��ٱ
��'t��� ��&����%�d�D��:f�u�3av���0��#�բ4�3v���@���,�	�x��d�M�aJe�#P!2�4���8��Xm��Z�d`H�u�� �a�0@�X��4Jւ��@�-��R�`0�R�  @"��G@I�cΩm���|��ћKŴ��d]�6kjV:,k��4����gw)8;��I��,c+K�9 �%��[�X�3Mؚ90�� ���Xk����;_$!��yڰ �7���!;	�jx�5�u��$"�$�[7ZH_*��c �Ͻ�}����N���[���-ڭ������љ����l~'�8�qV8$�t��1l%�)��@}$$s@o��|oF�c��I���F�I�%�y8b~p_��4�Q��!����K�VU�C� 	�%�8�����@��8x�L��t�JQ҃�";z��Z�dX�Z8p]��~��ɳSPJ+?D�����r��l�@�Ό�˅��-M���}�'DGg(�@b$���J+kJٵ���ߠ*��#���3��#-��q�N�&�D��k#-�I��p����D`0KBWv�d+���%����s&� #"�5�̗7sXl��ca�i���xn��k����7ZEb㫣�U�ݽ��h���uci
�/A͇S�4��ݕ!9M�9֑���H�-i���%�wv���xζ�!���b�s�f���N1�a�A�	�t�eV��Kv2�7]�Gf٤�^6�-��n�Vs9n��@��B�ܤp�k�"��b����Ϩ��m� c��H�a9#Ղ��؜�5�A#$�mXm�!4��
�J�OY7q��`�/��
���j�IK�cnv�݉):��eq7	5wTK��a,�m�2&�#�1�t��@�2��uz�ڰS��]Ihdݻ۷z˥���Ͱ��M�������C�q5E kj�Xb$4jz� I`wv��-�uf��#V�;P��+׈�4��v�+�y�U��8*m�!V��#(���F�	�ZH�ʎb����g8ʤw&�v���u�3��s�n>bM�)�H����ʚf�C�9���f���8�y�kZR0�n�YYB8Av��@��D˥e��x�)7�q��! a��d ���D� |Y�5�P�(���VVeĀA:��]d��@ړ�G�+4�<�H:u������K�v��ĈV[�m�m++6���	���� ���;�n�e�b<4�đj�kP%H ���7e�M[���",�#w\�f��1�8���u�7YC`1[�HEbB	v;��`%&�vr���iX#	�TDT1�e'��$"��\�) ��z��9Vu�W;RIV]ݻ4���q����Ma*��f�Dm c�)�t��є!�T��)äh��!��p	��l�6�1`A�밚FA�P,q^$r�Ab� 2��P�B!%R4#e��H�D�m��Km��;R��������;n���IK�훩@�I6�8C���I:tۓL�+�6��:�܌�I�H�"�4����)(���!�VBYBEH��F���ǭ,1�5����uҙ7F�2 u�X�����&���'v�%��!� �ġ��YD�].׶�&����4�J.$xh$��Qe�u+J��e�f�������5�FV��0�� ��m4��!�����PX'2�͎up,"D 1!8��%��&�\#[ ��R�;e�� ����XB��ќ3�#U8����i�YB.����!c���Z�4N�Ji�e��i��D�,Xe�ˑM/�Jd�c�&�ji���B0��d���ыickݸi���)���l#��D��P��Q�M׉L��Y�X�Ro�X���CD�R!8�G��bhv�m�ά�)J��[3QČ ���-� �&� �B&��&�$SX���l �@��LI�l1]m�1ZF M���N��ݥ��l�BU"�[��!!Lv��܎��a�H�+צ��*�cP�ìi/mkD�z���H�A}c��J��� ���(
N��k�D���$I���p��0
Ai^�f�n�m�Vp�tѫ֐ Y��%R1xILQ�זM5�)�uӌ� ��wWZRDGM��-�[�Q]#��\Z�ս���j�^� �\��C\DHN��Ȭ#�d�U�Y,�b�B[����wFV0������RD�	N%�p�M(M`@�	�!	H�m�!�i6�4ۻ��B+kZd�Dqۓu f�[lf����ơ�m�Ƣ��ٽ��q��5��:�2��� !���IG)[k����뉰�JB�9n���G������:�v�%��#۷6ia�U =P�؁b�iqZ��\���
R�QP��e��� �!n�����9������F�����8:���� �#��D�&�
��9ń�7i��!�T��r��v�)n�A���u�G4o�f�`qa�L�`+�f��Y��`/s�6h�m 2[͚N0�`�t��νN�&B�JG���iHM��)�D�#�����{Yr�.�.�d��i�X�a����.�h	�!V*�T�*�!�J Clg;h�ɥH���6�Gz�q�b�X��@t��A��o]���-��. EB9.��Qy�|u�g�Fj�������px �Y�Ys�^�� �k�e	հ���/k�HB��9����
i:�4�'$�IIr�����)L��c�&�i�ܣ� �$ ����VD�FR5�N$�j��)��{���ie�bJ�q6�Ȝt	�;q�]MhHHj���J�D�I���P���4�I��7)�ń'@X��tKk�����-�^��i���vͱ��Q�Uу���Y6��X��� ���4eR�XX2<ā�l�z�Zu�Ik(j����@��h�<�Vsa1gi�ԘC#�'�$6%F ��k"�뛬��8�d��&׉tXGv�Gl� +���^2��Dwk�8Չ����J@��.�$�4L)qM'�`:�(�"���v��ri�l�F �Y�i�M+�KT�qL�D\Ro2i7�BW*ۄ`����D�0C.�M!���m&�
�BUM��-�t� ���;g^Z�#�C�evά!��'#��i׻B�Q�8� ۤج%���f� NY)'V�� f�4@a�X��``L��L	���LR(9))	)��f1��G��4��1�h2�ݷkD�dI�5��۽+�HLv�&�"j�b �X�C�&��6 ӫ ��8�]`�%� ��1�B0�P�ax�/:&�ܱc4��g����`����X�Gli�P�6���M�����!B,{[���K
��!��%��e�f�D	L��f���B	�$��(l]&���(u����D^�2�F��ץmm�u�Y�4��#��.i{g]2����d���P�ǎ�8ͬ��Z�ݯ���M��͸��pہ`J8�YIVR�V0U0c ʇX��9�O&�J`֐�u�]�Na�"^���i@��H�7	5��0�a9��j�#X�;b5O�C�a�]l�YFB�^�Ba��8�D�!qζ�␨aѴr��w��Y���W��m˦'1�[(`�[K{fԷ#dULb��!���m5��]���ͻ�4 D�N:����  �#� $Q��	Q ��T8�;8�]�] K"EY# �TK DY�E
jT� s�/�yS�����~�O�|^Oq�X�Ǩ��h�}.G�VfO����h������5E�%!PQ�?����.1�R�9����Gћ���4����3i�*��!�EM-K���=����iz�>&n�w�p�0t�ú���d~$ϴ����P�6�`2����TE�\�ߍ��L��FS �t�Gީ�_Ja5Vs�ܭz@�_-qcU�h�=O5oe	�my6�u���`C�F��� 'nF ��@��AڬR�l8�����m�o�n�Ml��r	��"�'Bm��뛑䘆�^�u��m�O�^��7LGܱ�e���'x��oAG�r���"�7	�)��8�GT"�ED���MȒN[)3
g�l�s��kb�ķo�����2*ĝ����%YCh��Шbu�ѓ�ӆh1��[YY*��jB�h��Y�_��9(�V:�Lږ&�ih�8 �����?t�U��"�����y�F�Z��Z��4g��P�e��:"q�V�О)?�5���	��3�n�r�K@�Jm
�#�-���42ӥ� �'�[�֟쌺3�>6f���Š��֑)\J��}��i�� �a82���I�Dصa���[���L���e�� ��������G��\@Aned	A��aRCT��*�m��B��l/E��U; ,(��bHzo$S�ÍX������^Y�Zx�eʓM P��������'�k���p�*�ޅ������,v�jJJS�:S��U��� ��L}f�O�eRY&-uP:��������;��ל{0�t�<z2����S� ���{1lŐn[M;�MRt��$Y\�SN�+��,d�& �9%����c��C�QG5�ʘ�:E�#�������CT`��8'��̈́�*��s|p�nV�F{lh&j���C�|�&	���q
��DB;�,�l�y�s��є�B�1FN2�֒�~b˝�h���B{^vɶ6[�ȇ7!C`c�����9<���젶v\f⸒��,4ŭ�+�V�)�O�p5��v�5��PP�{,A��>GM@��']�8��mk�2�Vz5@����������K���f�h!r��B#��F���b@�h8--ټ2m��<qS�6Օ2	��E�~����J`|A:!ݙ���"���a��8,�:�FТ��P�S-�2�4)u�*=��[����$d9��b}F�h��n�,���ޛxI�t��!���A��;|�E�TkM�nB1��7�8�qͳ��SP:�p�̷#�pa��ؤÍ���S��H~�;p���|�7�ҋ+���1��bAh덖DP狜�q9�Q�a�n�yW<��=A-ϙ����n�#8pc���pڱ�Οr�7�]����C1i(���ga������⋂�!���(��J�Do.��C�H��4H�P�hx.Jӟ�A���ύ�,�^jXYC��b��V�����|j��eu.���[��~ű��m5��H ;`;r��X���u�^n�ۛm�����(��0�\��)��iR\��,KJ�,DBQ
��'C����s����t��+L쿿�៓���f<�a�qj�"��S�d�=��O�;a��c�㆐��������?�`�ؓߚ�D���f{�"Q����t>J�W+	1�����\A�O�?5�9���ڼzC��=��W9%�=�ɧ1n�]���#%y��4��D��f�(��!��M�rg_�L?����ZUT�����*(Y�`�U�E�݋�����	d�z��@�~�̡�X͍�5�C@��y9�0W�H��d6xTt���Ð8�b6凳}e����O��B����PϏ�0[ 9^Rh�����Fp������=���_3�$h�QR��L&�x���Œ�$q4����9.����f�&@�e�����J�:xo�v<��uof7߉-b�y�#t��	4]:����B�+��QoY�{�a�x��{�0w���V�@��>�<�n�U0�YH)�YR ���=L��$�ay�h2u���,]yx���%�A�M�f�j@���ά�����0})d�Y%K"�p�(v���	g�X�,!Ŝ�$�VgkA�r�<9#�ɸ(���O���;nt�ZpT"�!�?N���P��W�UK����N8v��X�I:ybG==*�g�^���FJ��q�u� �����#�5� �e�.y�L&��[�&"�йh�&Sy��\:�.}��B� pe��/
#��8]�O,�!�Q�\�ԊFIŸ���Di��{n��#�y~ $�M��@��1�3o��Q�4 -8�T��Sa
����AյQp����Îxt��s�� ��f�E@�A�1'��\5��ю��Y�҂���h�Þ`m��uc��P0�����Ѹ�a��0�D]�Fz�b&�lm�
���h�qM�i��e�Y�"���.vM@��@�" �٪������M�5ؑ�T���a�u'.F
�q�2��^!"��z ��%�f���f�, �j����a�	��C�p�NV2�I��vr�@��k�)����Fp�O��f �ڿI|)уƫpC1DS=<f�o4Ӣ�d�z�@Vkyi��2y��&��s�C{�D�k6�����am� ��b��")�nv�U��z�T�/�Ѹ�W�NI��;����Yn#}M>�!�2m�0Q~fu20`�G�V�`i���4u�v�"SkF,W#�T��y�=�Lɴ�����Z6Ӕ�oݴ���O����Xk�C�m�Re]����!�gJw���f�U�qE�BE��v��>5�3 �;�aZ���(��]|���������K�Ch�]����9��_�Z�"���xdG��!������
��KC���Vl|�G�y�ZP�B5���F�Ͽp
J	f;�������	�qH� ��8��:�ŇwQ�V}g�G���|�#�*1$"V�П :�W*�bE���%G<�� ��A���ݺ����3
�p����}�r�Q�R�4r�+/=�G��i �*z���rg�_~�=@�e�NBß9);��о	�m&�Ŗ���t�H+�x����,Vq�3Y�ZXN�����eI4r��+h�J4���� ���x(�aC-�ٚd9��_+��Ջ�4�*4D�<�)zoC�=�7��ۈ�o
ʳ/�sl��[m8X�����(v����GGW)���"u���T�_f[��z#���W1w�ł*��:n�.�6�8�×��"�%����Zs�By��@8M7(��M!la"��e!��Z]��㼖Pj�VDZ@�I� wA�z@�ATc��[0��ga����vٗ�1���vI>�*�*�G�	h�?P�2�KGlU���`�0�Y$�,n��s��)��˸�W��o..�4�&ʞ�_����2�����0&�U�0ޒ�
y�
�������̭���/<�b�IZ�sk�~�F�M�棕�)�5���Ѯmr�3u˵Κwb�C[nZ+��j&m�\��wuG"�\�nS#Sʷ�U[�j�歬��ҼT����m}���}�7��]�<��������)�x���ص��kS���-�TUR,/�� E ]JHUT 
�*0�� mP��q�"�"�z�k/� �hX�r�!B,@���������\�6C����ٹ00B��&�YL��8L���EUI$A���!5�Z���h�6�&��J����UBTaT.�@l�*�]D ĳ	�)*�Hp�]U!uTQ��d,]
�Pi`�LE��]A��)Z&���p`jb�"AP�����:+@�v�*%L�`!h)���(��:H\��/�Z�T�RD�)dF��Dm*	D�k]�@�̔
� ����d����J�#�ڇA�l� �(q���<(Ahr���K����*��YC?BJ�4Ⅽ!��D]E�@R\�P�@Śh-�W8��T�D�I9�!CPAGMB�1��#|q́��]�+�!A���ݠ�Mp���y5<�����{ 6 l��sQ���6.i��i����P����b�%�P��Mv���a��Z��E���0$*R���+*�*HM��m�Z*��h��#UJT��BhF�%��J(�D��JH�#b��(�ԑDD���Em[r�ZžZ��[��j��N�[����R��n]ݵmn�挖���6`����R �I�+V�j2����ǳɩ�b�e�lPO;�.�Z�y�^,YζX�&�[:��]��X�Q�cR*��T�%�ԫ�@�%����L��K�*�IT"�h���"T�UKQEU%F�R�A$��ATj*���5�n�QUlkk^+s$����TQ���XYoe�k[X��Gw�r�]�teDh�DA�$$2Z�*�� �ڭX�6SZ-��@�U ȷUZ(F-
��\��6"6m��۪��K�LQER�2F��u	PJ�J �`H(�[j�UkVR�y ����W+;j�kIVS��j浐�JJ�Rb�
�(�"2 *�""�ҐVD$n�[�,�\��2'���By�OmZ���Jې���Ԛ��H]	.�]E�$��P�Idd	T�P\qC� .R�tVLPB�	$\QP�[�/�j嶊�wVűV���o�TZ�ͨ�T#h�
����*�Ab�j�m�j�Z��mVUK�tQn� 6���e���Ǫ�+nU|771���6���r��Xۤj��j�І�x��t�gMd��`I�TG�b�c:�VWK]*粩6�i�\!am��<K�d�v���$��45D=^vRl&�۲����bBo;wjM����J�9|���K�ϓMWv�����mp) �y�S<���m�D �G�.�+5����׵�"k%���.f�	Vj�˷�q%'m�&�&n�` �k����ol�����w�������������w��L�+o�
斑���D���hKY|��'o{n�9͞�]&���	f�Χ^\gg!ƓF$!n��l!#{v[nk����u�r�����ԕ� Ux�`�G�����z `�p4wx���n�J�D�!���e&�\q�a;m!4�8���)4��A=Y�>�	��+�t5�a�������M��pE�}�<x�rz%\j�2i�3Q�!�T��4� "�<Re��p&�;l�`β���hq�n���	��D`��c��6V��;�9&��2���CU�ݭ֑Z/T N�8؂�R @��-,��*���*Os���'���%���y�2�$���']�3n�QiB!�Y�r�Gj���w5�FĔm[p5����:]ݖ�2]�\u�ݚn�i��a���V$�������,X*�3��d\l���h�+<�I8��T�v�1��H��G����[�Hѓ�#+-suM);[�6YqL�5�<�@[ 0��#c/���Dv�Ԛ��Qq�Er1-p!Q��n�Dsl�-3���m���f���e'6�1��g��6��uڈA�:�	��M�4�� ]��k�ڻS۾�@�-(V6%���pHG�$!W
Ș�Yf��a��'�rh��@9X5�ě�7m��n��-��u��!H[`P(k��LG�]9a5ΨJsݱQ!�����n��H����FU�WKD!�\Y8�w�t�<�0&%��Q AD��:����7t75slH�.�e�C���8�v��ca_�uꓜh� @4�TT8�"H"BVd��JOz�&cϖ"0u��$5��z�㴞�9�):u�'�9��&��y���M�_1�����yv<t�RZi��5p��G8d���Eea6��iK ��z�c  -���0*�q���H�&�١�Bi<]k)!�n�X�[��:g�J���6ޱ�%Δ�;{zv�[G��K+e���Q��B\%��<iy��Y�Ջ�xr��0SV
�6�c�a{���)k"�v�dv�n��ѪMtĖ���-@���hw3vR]�����Ђy����I�Z�$`��M饛�7g8�lem����t�����Rs������K�YZP��J&b@�II�V =B+j�^�؉�8�p޳m�la�۶Z!��n���6�!8I�ۣ�:oXtЀT��lv��8�K�жV]�Q "c�l%�Fʢ���u��"mg1k=doy�|j��LVgt�B۔^[T�&�,�T�`�6�-���,i�Q�,�eR�2+�Ҙ���)*D �����f��-���+��L뻡�@٣gk�i�I���Ƙ0��L�pT��. �L�Q� Q�<�*��F���Êg`�IJd�4�@̂�oS�ژJ�.��x��뻋��Q��p%6�H��e��kl��(%���B�lk�L�2��VZ �I���ṳk��-$��ҁP�X���s@����3f��m��6)���J�0�đ6�%^q|M�vZ;[!��Q��Ĕ�%�5��U�����a�����I S�tu���[a���v\pkCMljC���� JD,��0}Mr�&Ô�A�e��X���K1	4i���,�FT��a���BqH悐�Ylp�4D� ��WWVńIII���M'�WL��kH�cKj��jB0�kF�tT0P�#��ɸ]Қ2R��nG��F@��Ov���)���N�C��gn��цԒ�x�z�e��ヷn��a (��ѝ�cѯ2侶����u��ۺ	4n��tO�@	)h3G�r��H�mܗL��5�c#��m�������&�^@v�4���ڞ&�
�Q!�+\9su�-�M�P���%md���(����\�n�2�^,۶:R�wf��x{�a�������M6j�2�D�(Ul�c�X�%��}s6U�/������;9���=��B;z<��]�RNσ:��1����k�|+_
�z��N-�&8a-
�tdL*�Eo�-^����V�N�+�����
�7]BZH�m0�چ��t�@�)��~�Bo�#�`Qe��!�%�7�@_BlSI�k5�1��YeP+)�Di�}�~m��鬪j	P$Bd���nʙ��� B�{�ܟ�;����@�KI�����9�����}�]t$�-In�{o����G{�5|����o�p܀�����	��?ޟ[اuR޼�ͽ���0ڦ�)��@��t��P'M��G��� O9r{JQ�gЮ�AЀ�
��"9�� �|�[
T���@c0��� . 3�*nݩkg��?�@�?����;?���pֱ��w=�5Ns�&��ϣ_λ6#6����:�"pf��'�|�?�3���4E�/��d�b���n䰜��{p��S��\��)��G:�p�m%�~�>����/�V����Z׀9��8<���O�;E��Z�o�-��86�܇L11��Y����`�\mͮɼ��-��O�P��4Ѹ�2��i�itpË�R�H:h�Ⱥ�]��Y�?ZK�\�Z��u�_�K3K~P�����F�Ȥ�AJ��Lҳ��K�*2U�%����?]d2�}�l�b�| ��
06��Њ-�1r�j�-����[m��e�Y�4�Sh�X�cT�R����Mkk�j-�[U�kZܹ���o�~I���?��of��WJ�c�J�̢���0`7~g�0_+����������ae>~۷��_]w�⸾�֊>��D(,]ҥ�!"�+'>B�-� �PК���ׂ�v�5S5a5g��j6�V-Imymw-k�$�$L-��fW�gIc�����񄍺��4Pd�B���y�׉���&&#A���B&��^/f�B�:��B��/��nC��v��<k������!s�vΆ>i�f@��f5$Iu5�+�‵b����Z��o�źo�؉�[Ǎ^:V(�wvq�٪f3r��4h]�y$��܉�]�$��J$��o|�$���m�=v�����B}5��尾iK�h	|$��aD�GvJH��03b�bV2��+����z�S˭�w5�#S4FȒfE�ȋh�tĉ%&1wy��C��D�ηD6;��vޮx��jwr��E�km�m{���V�h�Ѩ�\�� �\r1x���U&M$O;��1�j�4�2y�]݄����$���Q�� $!!>c2]�!X��2؄�"s��sd��"�EF������* .���t����ҍ3wuF$��$��wD�<��,�S6+��Fخ�����}������څ����|���~��9���;����┲�a�_�������E��?-�χ��Тʻ�Zٟ���B*R�S���7ǜj��<2O���h#�?��c����ݞ���=��6I��"��d�N**�־/��ǪwW5CƯ[Ǫ��t�ׯ�I\�x4{�j&%)���κC��\B��A�D#R���m���qF@�HD��u��q:������.���<7�������l�'B�A��Y��{Qg{��Rk~Eo�w��C��<��\���-Cc|��2y��h	��*��s�?i�-;1oT}v���l��ߺ�x��rk8�|a��� #σ	I�=� v�A�����"����Cg p@0��������tI#�Fd9u��f"S& r�x��N뷝�w3@wr�$��u�2�D�B������1\���k����M[�x܋ƫ�G��r�rN���ci"f+�J&j4�L����y݌Hb�A!srު��6(� /` ^����N�7��={�{�*�w��̅�Rv7.ӓ]N��H��o}t�m����~�b��#�_p�<��u���?�Hz�k*K��t��/�'��%�����
9�n���H��yz��J�]��FJ1�5��?a��{�r?�)h�c�!)�1tm2��k��<R�a���J�%�?We�׿�dc4!֘�cW[Vt`�:�g�6h���Ze$�mӛ<��2����o�h��Z*�`�2�8	���>s ��R	e��F��Ԋ��G|o0����*���^*h�_]���Px�{5�TC���a\#s��RyΆjӯ���Fb�-E�s*���8Wx`��T)q�.�;w���ܦ��xMp.3�IKVYCko/�҂<��!7��� 5Oq6�����܂B�Et��D�8�}�M�S�Л�]hJ
�ެ/�-�lL��Ϛ�F@Ջ���G-ٟ�R�𙾞��E�9"���h~��A�"'���1!r��yy	4��ޜ$a~<�>|���J��5�8E��;���<��kJ��%�꧕��Tc�1'h��<%#?��G������ۓ�F��2���6M?�>~�(VX��UM�f�F��:��n{9Y;�äkVRV��:��
�}�O�۵�!{��Z�.�nak�53υU5�?ֶ�S�pf"�[��.ۯ�޹U�m	S����F(ѫ��Z%Ӫ�t��'��y�ڥ5s��]��W��	���X�#b��x�ga���@L�Du�@�y`�2��� �+�3H|-�Rҽ��#UH׬ku=�o��9�,8�Db�0��G1um����o���@�gۅ'u���-�}zّ�����'|������H�������z<��(�oU��!Zri}-�$�.����B��r��,�S�q	e��
�	u�M�&G��8{�<g�+��o
����|a�G��-�3`´;"��B�c3��ĥ�^K�Z|����X�fv�ő���Alw�ö��+�[��&'��DT4����Q�f1�>姼���_I��Qy�r3Aw�CqQ�O�NF�I��<��3�Ι'jE^��k�e��}a�/|��q�kѷhD�]Mae�C��KP��u������y]RnT��蔧uާ^G���7@��ZR����5�W	�PFǘE|::��n���bi����uQ~�'p�~a�q��rEª�;�z�hu�6$��!�
Ij�pʀ*�)	�_E��ίȤ���?H���Qp<��B��E���d�X�m�N5Z�BÍ��<��S���F.1븬��C�{�$U�n*��kv�9|뉫I��B������� D/����QT}}n��bV(%�ˡ=�<1Y�"��G�pL�q�J���p�|���<&z���LK2����Ӯ= �;	�6�Uz�j�2���,���)��;��9��V�ap�$y���UV�r�w�^I~��B$`\����q��p�1�M�Ӧ�{siiNG�#cO!<�2"9s���Q΢U[n��^)�u���Yy󘨤$��Q)c3Ѿ&���z�3{�oa�}��K���� զW#�Շ�|wT1�?�l,	W�}�9���I5�4�hy�[�R�L��׶H��Z��`�bߏ\�s��vƏê��5�_�~��Д�з��Z�QA���̙����g��L�F����� F�F��sU⹌Pb#�[����:�<�ء	��(_-�t�Iz5��������-��9�8R�Ѡ�0�Ԅ�L�ۤ���bN�i��^y�P��u�m�5�xܬZ�W6׋�6J6���]�z�u]���@��@)J����Ģ�e4�t��x�!�ux�5⻺L�'�˘��/�q(��Q��ּ[Ekx�WʩV�E�b�3BB�ݰ�A�wldLW����.1�Q�%�_.*,������>[ٴQ�1�j-�{�.m�m�U�Z��<$E1��0�(��M���x�$��y1'w�k�s�$�%�t�r�r�x׋�+�5�j6�(��j������3�	��c�X�"�B@��JH�
�Fwr4��Guƒ*5$jQ
!(�'Q�y~�w7��E�s���yO=�u~�zMqg~�O�~���U`�>�?����P��bm��-�G�J�7�z$�}��{��5��ӍM�Ui�fu� l�z� �i>5&��&��y��\PNz�4��<��zkVǋ���T�Qa0�::�c֊k	G�k�?]$�}��ސ:�����
�"P��P�ܳ,�w �ѻ3�<��~����M��!�ߪ���AOq@��*>T�V&����V�i����#��౦��2������Ѯ/�0׿D��b/5�ƭ��2�2��D���`��u��F���j%߬���L��u�L*^|�Ȳ�����%�# f��ܦ�� ��(c� ��u!�L$=G)
��OJ,���nS�
��x��0���e�TD����]Q�70��LCOq�(�"4B2	���,F"�A9��-�E��i\@b�P�]y�Ya�X�
)��WF*��F�MC����)�Je6Rz�wk}?;̣����s�r������ꢇ��u�h�0�d���`����u=�2\ņ7���f�U�9���G``�S()�?ۦ���C�"P� T�.���I<���Lg�lM(4S� @��E�S�O<��%�K*�p�����{o��͜�Ѓ"cE3lh�e��>��O��3��� ��?�+Q8�׷�QΞ���r>���.��������i�Y�|_+�Rs���3k�����DB�Q�G��}6�l)��e���ѻ,������ՕA���l�ցA�"��SB���jhc҇J��s`��c����P;�;�Ӓ	8����\��S9O
�qp�!t8�Y����YZƻO��2e��U0�V��J�yxjk��$x�6:�j�j�\��#DH�t(ďP���#�F���{�e<���"����Yf��K��皪F�2Ê}y�z<��:#��z����Ո\xr*��S������*�@�*8!3�_S⮬D?�-���Mz�P��w�(a@e_y�)dI�0X��X��e�)�>�u�ג�N���5�9m���я�f�9aZiG/�:e[#��

�m;������i�%�d�	U�D�\=�:S�^��+|T|}%�^HRZU�:�R˖2�:';3�?e��۹b�LZ��EP6$D1D	m���t�7��11&$�$�|u�Y��':D�
!\������X6K��K^J�����[ֹ�[\���x��Ca9q�� !!I��&$��c J1�A$��"-O;��-�h,��ȴU���(��~u�	��
4\�+����*��C�ܹi/�਌��Ȩ��µ�j�J�@Fd{�z�&�r�Es\Mo�(�-$Qr���;slN��z�������[q�H�EF����/z�ш4l���ƼfQT}�\���F�-��=���R(s�'7DӸ�5�E�w���r�+���j60�|����kx�:-_=��N�q
ɍ]��QlZ�FƣW�������Q��p��QTlIh������*|v���^6ܾ>{^+���"5z���m\����VD�Dj(�E��ѵ��Z������E��oA��H�\�mz�m^(�m�U�1`�Rm���Q�ޢ5�m�+���j��(�ھf��^/�\�����4�)�O��#�S �&o��ŵ�N�:�Tj�\���ۚ�V�ߌڷ�����b���0E�Ƃ��I�hH��X��snW~�y1˒�2�sq�Q�Y
*�vᣗ4L�EQ�d�Q����^u��t�8J ��(�KM&K@XƄ#AF�!�mˑa
O���U��ۚ6ܙP
P��Z�KEA,Da(�ʤ��t��w)͒7'v�ѸWnu�QF���&ww']3]�ù�C��k��]�]���5r��NRm�����Ũ��uݵ���\,��e�i5۝ҧnjuՇ]���ۑ��ff@��221���t��;p��:!lA�����W�|.Z(��F�m���'�Io�j��ڞ���1Tj�=�y6��A��s�Z�h��ljJ�s[կ}�,W�\�6�Er�Ux�E|w%�oU�n�� �A����T^-|��j�[r-�®�:�Q��Z܊����U�|��UE�xx�񍈟Gcsl�/�r����hص��'-��5�����u��`���bX��+��W�b�~��U�j�{����!h�KU!! �8�Z*T_�ѽ��YpWC$�EΙ�K��	d3 �-- ����͛�j�?��z��13��J��j"�DR�HZ5d�[������ZUSQ�dA$�	 Y��f���j�/�k�6��U�6��FK�qM�y�W����Q�D�5��E�����{��J�ӱ�^s���w}*Ǚ�7?��3M��V �$��$2�Q���j�2wm\�T�"H�� �:�@���M�wI�����k� ̀gE	T�n"��
�=N蓻�Uc\�66�Qb���G���Dd�	$[�߻�vf�H��GN6�U��K@K�8	o]���$i��qʊ43�9ͷ˅Q�������/����o��7����s�1����P8!�
���mo���b�I�JA⹣L��{U��fđ%�Q��n5��b�Z�}��筲�gg������F"�04�	P�Y}�Z���^��m�s���r�t�2����McF�E�EIY��"�� 2+ �Q��9�����c��d2c���'�Ϲ���R*H�""	C��jV�*,�	ۻ��7:��}�e��\��⹄@*�D$�J��p���N?�ۄ��5�u�xӕJȦ�P���v��k�{���-��͋r�.nU�t�Uٚ`�B�Q7w��j-��*,TH�����;=[rWn�����F���NC���l��n��_�g�E�"���	��F�Hm��m͹�إ$�(�cA�
����F�%E����UxՋna�g�/ᴾ����	���3c��DP0��$e��*�~��P5�@�j�(�,֍��o{��ˑ�`��V.%;������q�8�wǛ�����t�s�E
�?�}6����o�u������N5D7 3�uW�׊�ѮW6�Rbf�9�b�/K���^u�L��A�@��h�9FغZ�UW%�m�j�Ih�'�l��Ǖĩ�!"��J>��k�6�[^7�+�Y4Y��"e��s�����!C^wI	su�4I���mQ���k_v��\ QD"�B��@d��m�r��:Q��U��\�\��n\�0�u�1<s��Ji)���[��W/�ƫ�Z׍�_�E�4��|��jjA&lh75͋���$&�ǯ<���t�nG��o"�wK����h��uDZ��-R��H�@Z��Z���E�N�G�EN��x�2�"�p�1��0�!�ww\N����(es�l Ld.��T��т�U���m���W�&��m�^"<U�ŹnW.j71��v�ˈ���& ·��=��1(�f��bb� �w\�l�G��)qIP$FE$P�n��U�r��V�mʠ��r�h�w�h�⨮k��3�3�Q�{�c8B��N�Ț`�"1(0\�4LH��rCJoWD��E��o������R���H1 �[�%I/��d���k0%$�2*02S4\�[ˆw$�X�7K�!$N�l�v��Q�=�x�ۚL�%(�P���o^�*ǫ�k_�W��KYAU�޶�ۑsk��HV,1� �1UBs�4@�j
��]"3��wvXD�1��@���+��s�E�y��q%� �~.���5c���
hyWվyH��$bȬ�&4�
e+�i����m{f��m)����M-�b:b�0�	*R̓$���BI ��_:��r�x�S6��J�����~g��?�_���㼷�}���|����|o��K'��C�����@?������e���=���}��������<?��}�ʟG�_���y�q\�ŗ�A���l\`����Z�$N�� L)2�J ��т!n��qs3Jɛ���"��������DB0�L�t�礜�\��8B5�k���(�Cr�e^�^J��i�*��N6�΃p�J�:L���n�y@���O�hۓgd@�B ~huwl��v�m}��S@�����T3=]�����s3=�~��g�g9��.��n�g�)���i|O�?��/�g���"k��l�:k�������ln�� �{��=�Uos�5<�a��_��g�.�]NNo��9�[���^k��r�f�OK�ou7��/�S�#��u�K�R�����������WW�b/�^�~���[��e����t�7�/�p��;�g�  �i����L��9�f_O�̐Ђ��g���e\���ESښ��J'�hu׳>ޏ|O��L)�$�ؖ�<��=��G�}WT�z�=�S,�hx_TR*�e	�r��b#�BT�/��tD���aW]˱I̱W��6��(�G�ς���=���~��A���_j�l�N����E}G�us���i�ｾ�ƙ�~������7`_�9�x���h�y?�(*�{��f9+�W��e���T���=�>����i�[+ 6���N�}>��;�f�*JT���	@���N�Z�mN cO�yWX?~r��a��yRK_�y7<]5C�;�U�4.��Y��Mso^��!���4Û
#2]�b}�]}�h�����9��%�D�mi=����1Q����Լ���R=�/MZ�E��% (��Q��>�:Ǽ��G�vL!�&���NqU헛;�nМ�ٙ�� ��=Tf�eL\�$��W�pq�a+\�:v��y��l2��gT�����%f�o� �C݆���%}��oQ�m
��;y�C�n_��Fކ�QQ�A��/���V���3M��zf�iS��r���%���,4C��zyc؝NzELW��4-��I����a#�%�a3��ߍ����3�ߺ�K�r�V0b�u
����j,�v�\$���̔sdW��2O�t~��0)��5I��?;�qw��}��սM���<�8e�,$��A��������5�T6�&F[5���i���:�ɟJ��m6c��\�qFa|�kR91�S�u#L���<����� ��3��߭����_����c�%,)���!�v��p=���D����O��(pGv��ع��P4�t�8d�\�t�eE2<��{�-<�D@�]r.�>$�iA�P��3Ї81SJ���O�~!h�*x�H�w#}-��O}&�	#��Aټ�t6l(��F;���͈��qk��'�a�q�����	��a-�+"�IvCz�G�����?6�S��T�����!�2�yz!�%��]�b�ӻ=`�����X�9;����%��t��[V� 2�'�ʴR��a;_H��g���٦�1��Y��'�0��;uT��)S�B��er�Uq�
H0�4[�:�TY������7`���=dO�e�5f=d!���XSfG� dq+{:3�z$��@�v�w6��\cl�uņy�J����d��h��H`�/�������44.��S��^򀩑�r���&�W2�,c�(�m�$�GoS��:	�'�E1^�9ؔ��pП�=�*m�tO'v%R7c�+�s��.����K���iƐO�( �i�Wvr�k�7�k�Ŝ�� ��Ř_�1ap��b�3-̓�?n<��D�{9�Ϧ���*�3���(���'X�����̥5-����Q��x�2_H�C�޸�v�x��P�'��Gp/߸k�_=��ԯ�MH
�8x�i��Y��K�����(�?]�ԋ�2�Y��<��P����Z�����V��V���䌩��&�hD
�~H��2�j]�I�� �O����hL�l<�=u.�]�Ff�K�Е=���=n������M	_�C43���
�c�?Be[^G�Ŕ��ћ�ի�Į��B[���*����z.Y�'�˼lq��A 3�vq��@+ѧ���v��}n�K��,�5Cٛ��2�K�H��%�u�T���\�%x#���ZG�ю
l]փ�� 7$��&b%��1Bxp,��×�#~8z@D��������+<�@�TE�nj�m��%�| ������C� ��� 1��5{�1W���@F@RE�����z������\��7���˿��N�G�����q,�m�[g/�+���a�)	��'#��������.�b;p�����6����yy��6������wm:z~�×`8|�n{�Ǻ����C�X�}{��Q��'�ǂGd�$
?���r����R%R&!S������И4����Hthp��<�g���?��p���G�P��q߈�I�:?�����i�8��ۗ+��:p�ɉ3��>-���%��Vϒ��{��>���r���Y�fBS�[��"0H�p�( �0�rˇ�l
H<n̒�R�h���!#`�T��%ĵ��M��1��!�����i`h��/���;�[��4;���v��{��{�� �8%�^۔��R�
w_TRu��1�.��x��T�`&	�J(I>�� b@Ҁ8F���KQ�'Z@�1@�[p����H�bɆ8�<+�Ў�Q.�a�K���
N�w_Q%i[��XQ�����n�GF3Zj���dFэ���E�AE8�W	����oˌo�z�o���}s�	��I��}�4��`T6��g����mF_��;����c1�|._oያ�
x���IK`�W�k�>lʦ,Ѝ	犮��ؒ�Ê�����T�|
\\�1��Ղ�R�n%6܃��mͨ?3�Lţ* �L��+�Gç����lMb��EF�J0L�����{�(�Ȳ�be݂��K7�B!G2Q�2�z��1X�˚��ڡ�`E�r�����O�\�x���N��fh%ʎ��4.M��@��ڭm-n 1+v��xԀ��$Q�`f�5�H�,œѼ4���P�-��^$�E	�MTevi��a�GSi�m����A+݇uLn��X.��!�W�1� Rq. ��/M���_��e����i��m�MU��_���wh�82$����?f����"���}�f�Z��;L��k�=l�k�$eEP�"t ;V �J���B�$�%l�$)� ��ɓ��8��"���*�E��;��V�X��V-�Z�l��c��N��˴�������?O��n��y� \^V�}v}�M?!���S[��6W�� ��xo�.�y��(����YR�΃4�o�߱O�F�i���Gӛi㶷*���#���u��|?ɽ���c���L?�'b߻�˧V1�KFm��<LC�~�Ā�*FHĂ<hBH�fʙ���MO���!M�$	��20�H v�
��l?�麞�}#�yM��[����K����g)��N���o��zN���Q�O�+��u�a�iaiU������׫}Io�Wn�32�$ ֵ�ks[�j5mbֱ�Z5�*�cm�6Ѳ��B��� �D��b�	C?��o��}�k�Y6����m���}_���[�r�G��|��|���o��P��W�Lؚ����6S�EߝV�X%d��	����sVn�%���C��o�����{5�����t�����x~��p�mu�:�D��M�S��ݫ��+�..~�ٰ_<ێ�v�E���l>���v�����eJ��A�)�*�>�s�6J,T��l�G`�+&yv�*���x����P�Խ,�� =�ˢ�c+�V��Eu\:�үI��,Oy>W.���Qir���{w��ޔ���I��G�.i4��--N�8Мu�����/#��A{�P��bb**#{j���k�{;%�B+�:r�,̍��kNBY���E_Rs�L#K��2�_"8��a6��6�[&�,e+b�2h�kf'�#��3���hI��)]��K!:$��铻.��V�U�MR}{p�Hx��T��+��ޜR����l���0�����:@1�ܙ}�-���i�X���׷�t�Ԟ=�zq�N5At�{a0���N+zp��]�� �'�N���<��}H�}4���v���԰v�X��x�&���w�������eC�b��z8��c�*TU��٭�mOi�C�=6?����*�s���*C�{|{ ><*Ǖ�X��$:	sh�5Z/W���E�&,Q*dO#a�(NoL�=u�k"�`Dr�yh�;�yԣ(9y�Mw��al�ɕHǗ���T��b�m�S�5�}�SqՋ���3�����Ɂ�'*Vf4��bk�d0�FQ�jĐFl��,n{!�a�\��w,s�Q���o����Ŏps�K��ʶ�N2aC���Ԅ7GC�Q�Ǩ�������s'
W,J`U�E<;��[�0*��y��fڑA��{[3�-����Y뀡�o�]���.��X�a���gm��~Ó�[��� Ø�`�COwtZ�`2E�HM�^�o'ɰsZuwg ��2��NI[��LH��-��h���C3�j[+N��xs����Ik���I-S_<����G����K �~�qŭ��]A�wQ|8��6h�<�
8�q���G�$�a���ogZ~>�T.�T�ۚưʺn]4W}��z���&'��R
�C�����j�Toe��j�4��T�ϟ��"+�/��B�K���m�.�p�U���d����iJY���#�Y�"(�����NT��^su<�|U��j̡��*A���C~�$�]h�Bcw��s��Z(�}�ߣF\6gl��{pOI|��l���#Й�?S�TIuB����-tS���2v��	����
��م۸�s��UJ�0ݠ����]X�ٟ�@���2Y�\ފݏc�ꄄ#�Y�)�.$p4υp�pP�R��<�؞�6m�_�-�q��v�G��G��-
Ǌ�okIy�"��S�ߊfa��N� ��|�N����Є����?\�GD�-��绶��'E�x�r���q�m{�/��F��tE{udO"Λ���u��,P�':o���'�G�ʹ>v��i}+��|�B�5�D�
� =�:&@}Q��\�Ω^o���Q�$���8����Gc��Xrϟ��b�J융��u7�3��0�[���;C=���Y�t��m�;z�.�};e���P|�a�E�Q.����x� �
�:��S`��<�gM�a���U,N�f�G'�e�v?�V��I�-M�ؒ�.^����#9�^��Ϟ$���3ӭL��k)ww�y��S�Fcͅ�r}q�{N?]�+��0U�&�
5 xSD��h4t7�F�]���<�G���k�~]�)��~gi��6�v�D�Dr<��[�B�nmm-��X$$�����J�B^俭�+�^��l��|�{�7��m�x�ܠ��!������)\t�7F?�s���s�����I%�����oҧؖ�?�;�UD_ԏ�YQ��>C�nX	���.��J��?��e���8��4�%�~��8]��P�����`̤�M=`P�Qs���16���?2�$��)��(�?����`C�A�r�*� �݃�K�{eC�Ѐ�<KH��YA*� T��Қ-Cm�Yt��N�`ٚA36db��C��w��n0�TR�`q"5�¦�v�&3�\���B㥒�0]�*���pF�A�}1n󢼄���}�/�c�Y��������̰#0��,E�m�xZܾ�{�w������p�Y{W�,�=����XQ��o�Xm�(8���)c�,n�	�\�@�@	��X#���Sz4�!���Ĳθ�7ښd�{����}����*#( Pj�,�{!�!6�J���	ڵ��\��_}烖�
{b!y����_�rv�������ы綿f�~W�����O��1�4X�9x�{a������>Y�-?��[��Ј��[8�9�\�}!��s�<Cr�#�Î6��Ĝ�E�e%^�Yb�戎W5��He�lp�F0�N߾��w�nb�gή�>�h��Mv�|J�7������rDl=��R�XY�{G19��n�<1�����b��ĸks16a�QF�L� �ק�1�åp\YY4<d2��q�c�*�e=�
V3�X�1�8�"�4hQ��Fe"�1G���\�,�2��aH9�d�� 9��7�y��"5����b�Y��"�h��t
u��i�P��?%E��dA��QT�	j	���jy�]�]�ncG��Y��i�E��ĩ �#�j\������%ΊNĸ���d�ēؗ����2�b ���(��d 8eAQ��`D$����}�F-R��Uh6	�dJ�^E�*'��8���_�;�}�ӟ�=W��>�/y��_	�y>��sG��繂��o����.�Tvh�	 �2A"(��� �(���ʐ+D��`�D ��ovO������>��|_��������~%Y|����rs�����J��~`_C��������^S�c������oO��EhkoO�𻙯�����8�����v�񍆠���*Q7�Y|3e��� �u�����@?EQ��o��M�����0�)����j����1�u ߤB~ �'C�
�j�y����K�Hk��/�����w���u�_Â����kr����"��X�����Ӈ�{-�k����p��׍�m�����������M�άގ���{No>�v��X�*4!��EZ�/g,ti\F�6}�T9>Z	-$:a��؈��t	ba����3@���·�Ok��E���k	|�_�w����)�-�J����Y��Ւ�<�z�cBL�H�n>��Sh"2�MxQCg��Yퟤ{�f�Q���@;�*"�#.��)Y���68ƴ��m�sŭ�8�̛m�~x7��] V�B =t9Hz�;E���	�~����ȇf1*�VI�I
��a��17st�;�>�e��O>�[N�Uk1�v�zM�؞	:�,�uzh����"����*�Xn�W�_Hљo����b4,����O J��Ap�]^d�L&��� ��'TR���"#���bu��i��S��>jl���Gu;	�L��,4=�r������m���rj�k�T�z��:�S�|�#e�=v�/��ts����R�|5��ub<�Q$(���5��"���7�M��E�_
9�ӷф�.��4��Y\ڭ�.���j�9u��r��O��9�X��pV�E�e�s��Ű�,�ϧ�k���R��E�mB!�x��و��F�#[	��=�!�����Q��A݃2��:k�؞�0C�æN@���P��2f�"H����Ю��5]"��M�*�^���KK\I�b��m��r���\�7T����SÎ�k��"/bfk}���DVQ1@t�������8Fy�<´J��ύ������L�"5���ts.�q���s��U}�\���ʄ	��3F+�ξ�n�)>��w��!��+~�a��o1LMR���%x��� �v��r<�[;T����@��jH�#1ExRy�vL�+���~�/L��E�v5��	���%���z*�ׇ��#��Y� љ��y�!Eýa"�3�-J,�N�w; ����@�v�OX�B���[�-0��@��G��0_����ЉM�v��h"�.���s��I;��x�(zWS3������5�D��;B�|t�O�����,+"����w��uܖ^�;[S�bY�xȇ bi�Mc�OR��4�<ۺ\i�ޥMU�y~]�}aΦR_}w�T���j&Md�ܻU{������1��?Q��"c	���kw������shB"�E���=8ͧ���y���M�3Į�FBD'�ޭ��P�;�Y�$�.Gu�.�=(Ǐ��A&1�������5���'�7T�`H�J���-�%�\J�҄
Xw&������O:b*�??Q�q��/J��a�m��n��9��C�Q=eaT�D�"�.#(�BvA�>|�#�z��XLy)�i�7))MG6���T�*�R�qƛ�.�)rT����L���zt3�]��)�N��d�Yhm�-~|��0��$����:���%@�a��\Z��nw��N�ʅ���^SS{�û��!�c��;y=�;�ĉ��{ψh��%�(��jW3{��b��E���d҇�u���Z��UZi��}a�V��^WG�z/fPD��mBЅ��zF��r>U���W�=\~��j�.[��q��{����e�-�:N�v>:(t �g͗���o�T��2���sԢ���� =���e��i[J�l�*V��� �����u��w߇�@��d���p#�X���>Ȏ 蠒��;?�rw��"����ԥ��6�������r��v�]j��>m�=��Q.%nW��˦��8x�4�����o=��-��]��ӱt0�8�W��*��k~�'���s��zy9��Qt7�z($�_���S\s��,�l8�n�N�Lݳ���:'Yh�Ɂ�B���ȏg�m�
�����nw�����)�*%�eDNX�C2DF�R�b�T���X�K���|$�}s^���f��뤽�B�԰ei�"xEH���0[���=-0�d�㮊�2f�!��j�&d�U�5��	��67T<�eyW�	�eV�ڕG�i��`P4��Q#��>t�SXA������0����b?y(���!?�M�o�zɲ�}�u)��R9��F�_��Dr���4�c[7��֝>N����=��������%������N?^\��!��m�l�Z�^=�gH�ة�K	�3-:B2�²z�Hן]@0!�}u��,�<;7.�߅7ٳ�S�Q��$���׻�ǯ(G�wk9Z����uqeYj��&������o�+�F��|����	����/9�=-�����a&�~��M��Q����Y$�8n%�~���t~��&;}��|�V<y���`����f�w~��*��Z��MI�nu�m$�����BWj������/2�ŗQ;���*-�(F::����8	,�>rTA��2�0�|��H� ȶk�n��<��=�����C:�	����~hM+�w������l�M��1$�A*$�!��6�Rk_{m]$��yt��ͪ�f���Y��;�?��Q����\����3�{����r'���I��~ߣ�3��N�ۿ��t�7��_#�w�[���Q|�Ǩ:C�B���No�x����N���7�t7�!�O��y�G����ޯ��|�/�&�N1�����{Ѻ~�F�-n�� �5���H��,�x ��w��_p��}OĳC��|���B6�� ��w����U}nҡE���ڟ~�CY[�P��+����PH٘��QK]����l
���ܟ�k�~m���I�n0R���z|\�0 ��o`-<s�6������8AL6�:u	�Y����_1��~�QCx�ʀ����)}{��b��"}{�y���
d
nX�:ۚ��a�r�p��y聑5Tq�b�����?n�n��{�ȫD�
:[<Kڂ2�)�j{��@�����ڴl#ɓd�J{���V�;Jٹ1��n��ܪ���jD8��Z
R�
���bt�=3.B�^k vT��%�l]G�T���w��:<�u�WB��_�=.	C�Gg�c
�M�2n��YW�DIg	��M{V��@��fǐͣ��ӳ�#���
��ݩzMN�*ף��h6@��Ĝ��$���E�����U:�#�>��$`��8���a��N$a֍R1�6���mq���D�OjX�՞Bu!!z&�T��
�4L��o�K��i|R�FC��>�p�J���݇�"�}.u8ڀ�4g�;���=yb���:j��(��J���U�"�BN��k<`I#�-���"�Y�/O�m�o���!/ѿX�xr�k���}�l��
B�0u�!s��Y/�zP︩�5Q�B�pÙ��� ��k��x�\��#��!������CW���C'���I�l�+��L�)�Ck���B�J�*� ����>�������+l��^��Xebn�Ħ�ZRb
��/�i�ڥ��Cl�ug_�g�?�	d��T4ov�
��N!��+c���0%am��[�0��w�q�Y�1�k�^��8-Ҩ�S�͘�-�>׏��^3�#�C���w�凓�g�ׯ�2�;b���p[�O
�ʣ������h��5�d�5c���hU�c�Pr-DXXs;b�쵍x��Ot �sL^k�1��ފx��֢/�	w<�'��^�c!x�·5��|�D����M�>}(e� �������h;���IZ2�@'w5�
f:T�u��Ӑ���`~ޯG�T
A&u�Kэ0Yil�XF�u*�M��G��%>�v芗L²t�Bmy1����
f��;A�fV�͸x���l�T��މ~��j^�ȊrE�}���&AL���J�ڑs����"�]r�΍���n��6�=�աwu�f�3sx3:oM+�p�7���W�CR	P�#�t~�Ǽ�ؽY�by���j�sIK�`�z����O�P)����׮�m~�$bbF��k��6|?�v�Ɨ#9|AG{�Q�T]��6�Μu��`��iS���"d�J����Y�=5����\�CF�6�b<,�wq�*�<�R=qê�-�8N�#�.�՟,
E�L�*-0�J�e�-���+�#����b��H1�`����L����W��^ �Fy���`��f0+���E_<yNwdBd�M�h��d�?C�c)�E��&1]]��VN���1��p�^�]"�Q�c���IbW�VӜ�}a�>�wO���E�*�8F�
����-L�X�[���1��Q���Qfv�L�JT�$;�_w�`ֱ����'�Av-f�hD��U���I��tf�\:����c%���G�;��4.rXBҐ�'�?����Y�ֈ"�6�ht&��S��G{M���%�)խɼ��rTl/�xɿwU���  �{4��������W���}�7���;���C����IX��iw��&?���V��2�~|?�L��u�-8o��˿v�q� ��O��i���o�hǰ���avQA�r��4��Qd8p�n����g'���������ӷ�kLv��m�a�C����Wտ��n;a�ۿ=7����Lo1��h��"�H��s��h:^G�;v�v홴'���O��@i2�n�"��b�N9tx���B������TB1Z��kR��##���[�eI���t���T��zS�j�(�D^�M=<�S��~��_����&���8]�z��c��q����l�x��0�w���	�z�uza��ٿ�M8i�׾�{qϑ�7�*�O�R�IE^U�8�H�
µ.��8��������r���9�=>�����_���*��}���r��>����r~i��~�Ma��}_Y-�V���.)�.y�r,� �$ �T�"9ӄ��u
i��_��� @I�QRo�)A@잚�1�T�&�tH�L�8��X��Cp�Q�uj�O�Ѵ29|���~�/.xvk,}<n1�/�}u��t��ߞ<o�'wPRXU���#��/O�^9�O�ydy��ۿ�U~�ڨ�����	SΞ�:x�� ���q�1YAB��i��U���mg��v�'p�>u�a۝/������Xuێ?4NO��n�|k�Zw��h�s�����vX�H?H}O��4����������n��>��~�����߱}���Cۯ<~a����cj�	���5v�j֥l�b�2.�P�Ac��,���"���#�{~��l����\>��6N���7�����/��9.�����?�>+�������w��=�����w!�ۊ����.3h]��dÌ���3O"Uм�������[­�Eظ�Mʚ���-n����C��R:�M�\��!�����2�NFT��"�ga9��յ�I^��פ����J�d��t��5���E��݅n����.v���4c�1�q℩
7�ܗIs�VT����Z�4�uWUQʡ�@�c=2	iL.�up��Ԯ��r��"�泻Y��a�0��m���"���u���'�pB(.�6��D�;6� :�X��C5�/:%n��%��tL�c���N:�w/737�����v�eOe5ei�[��/D���u��(��"��#���t�DY�����#�Q�n$N���WnC�rB�O^��=�e32�9�>a=�Jw��a����ˑ2���*�
���yb��#��`�W�\���x�����	WTH���]�(L�+�ӗٕ׽�p�q��v���ƾq#z�o��e,��L���cP�y�{��*���br�n���}��5qZ���3�d3<	�#a1�P#D��]��s�܇7�_G�8��t^C�A���C�'��
}���"M��w���D%����M���=ύϋ�~�~��fS���8��w���k���SO����'���)�K�b� {=�17����Э5��v����g{Lo}h�J0�$���g�[�0��dE/���F�W�_� 4锽aX֟�_��&�y9�=���/�3$�{�în�r^e�t\��Ч��UKiR��Q��	Q_	��J��� ����A�w�[7�fr��h'8��;6��� �ϩW�ӭ�U�v��A;�:�3!��{���m�G�{t�;i���ּK�&�	���i:շ{�A6�N��%�4��=���y�9"�Ǝ#T�Rp���|�������?�cup�O=�����B8%�%�C��u��mZ�a��*����������M.�WuM��a��<�C�s�#H	��l��	��8Tr�!����J�˖���}َN�-֠����á�,����"����l�V1ϟ���`yJ!�wc��9���Gݺ=��q�yv���"�-�5>�O�i��P����=tn��\B�`�{	>O9��3g��D��f�	��S4�.7`�,C'��M濽lF��
l��uy� ���L�&G�S@c	�^C{���7����7�,ֱ:fb��OV)@��0wV���
�Ԍ�bz�^�z?`ֹQs�yZ��V���vh�� �6q�+j�\��x%��� ���C�1h�üz)��^S8�����=�o�t4#�dA�T�S�1jjf'�~�-χ�j]�=��w^�F��*��H5�gN);�Ӛ!�A���M�«3bHc����t:0�4��t����/'�Q]��<�}x������Z��>���ߧ����S1��w�u�<u�/mߣ{�\��N�)"lDU�mπ�$ib9��a��K��̻J�ש�!9��J��q'�'�|��v�%N�>g�P���?]��`�=�]���GgP��ø���&�Fą��RB��B���{��Tv���HD���7 �7�d�7���8�ԙL���_�{����&�N��۷��i�u��I
���/w{퐯�X<�U˾���;�C��v~�+�!ֻ�	��:�3#��f'�X�AP�b6i6K	���z�s��3t���Y�� ��'B~UE�>8��"��m	;yz�u����w��zV�MN~}��fF�2S\�A�!ۘ�{�#�Y���{�0�����BY$W��Y���A��L���N�ImTA�Y�0����^۵J����� 
=�9�[���o�a6 o%�ʮ��a�i�T4-������r�v]�[�8�����~�$���u_C[�4D�&r����ggj�m��W��/�z$�}WGv�v�T%Uo�#q�4����ɖМ�YJ�iw��p� �&��F��Q����@J�F����|�{e��{�k����qw0�:�Y��QE#X[�3m��-V2951�fbWd��/=�;c䭮ߢ�4}fCxh�5I{�S!}�R��qy�$.��	��øP �.#��t�O)�Qg�8 �.���Ҹg�ߵ�&�a4Y������Z+�SHiB��c��pRT��B�BL�&�՚�֑b�w��ObtK`��XH_+����4���ړA9 ��u&�]	'��iS�*�F'�6��f�@P�j�JhF�"����fn�(�:�U�y��Itd�<D��='P�]����\zn�^G	(�e/t�K9��N�w��G�|H�L�0�+�Ol
 ��A�y�4�xf'4r7t e��(��~�uD�k+���e"d����gv˥ql9'���:���H������<�H�F)�Rn�{A�� ρ�_��?��`�����eIqxC/׻���W����A�{�}X�����p�]�x�\��%3��s��x`���%���v}v2��Mo������#���|#�p�l���������+��*����wMu��Hv��8X4������u��V��f|�o�q��k�\�N]��Pt#���(,��ۿ�8)�?'o��)SA�i��'�����7�����a��}�d����{�����j)���K�I{��0�t��X��d�9�:��J,�q��d���i�%����Y�z���r�ӝv�e�|¯Hq�
$�W��['"��� �� 	�u��E�M��k�1���L�����0~��oӝ0���������p-r������o�g7���ݜ�j$e9Z>^���cL��Gh�K��'1;��t{��	k�S�zq��+t咦���s%���{���r�|=N|tM�/oO^��~��,}�q�t���^�ׯ~,�dz����Q�������'wO�u �vY��
�Rh�ul��Ǝ)�˗�'�]^�/i>֏���1GV�8|�����O���֟�#�������ґm:P%t���}�ǧ����l���y�Y%Z���V��~]�l����<�Y'�:�n������,�d'����p��ط*���yd�/V�Wژݣ(�*�{eߧ�D�}���o�6�u�;���li��Cd�v=� �6H�X��b�@��lhn��� 2Q��-��+EQ^/��紶����5��@P��z��ݺ_w�|L��|�3��<���!�?��?=���W��{�����I'�ߕN~ݼ���p���]j��Wmy�ݱQO*��YV�1Dh�1�&"�r�cŵP+)w%b�jq�pu�E˚����xb���D�
���3��#ccMEh��`����.�������J�:3�TM���s�X�V���b�9�2#+�{oG	�������n���v���j�\@}��mu��4��W.��f�jY���wk�-�[����3.�DLT�+��&ݬ�c5��y*/�F�zh�7�q-)Î���x^�6�es^=7+/�u��r��U]�[��k���52�F��G0G
�҉5R�I�U�U�Ù�cc��U[��3��6����z�pWO]�v�\��sy��v+�oEfJ�|!,ʬ�6�w����05��i��w�Υ�b��.��b��$��e�p�z�]ɣ�:`\8��d�و�'d��7]JU8��b+:Z�=Ź�#F�jH�Ag�mK�<�U�u��V��52v��TU2N�0�r��������ך�N��.�UʢmT�]��q�iaJ
F��r3'�^p�����5b0����㗓��&^1�qY�Ҽ�geK��k�y1�j�VdvK[M°9br`���6�7qt!L��p9Q=Qw��|ݞ2���K�j㻼�U���(j�9p$a��k(�ˋu�Z��%�®nj%��wY�X/�)�)mX���ħ1Mk����gY���Tf�]fI���w�9qEwT���o�ff����Ed�ѓ}s<��'#�`���{.Rx��0*�uSc�,���s) �ۅ C�	v��
跞�x�S��|��x���t<�C������6^�x���x}v=w9�5�~���/-����=�T���O���?7��~�gK,��
;�Ҽ�����}�xfØ����Y'�7�j�`������/��L֋W҅�=QF��M���5P��}s�HK������{�_,6�B/���Z7�Y�"l-�����0�B��kd����n�nf]���T�G�/4�@%��;4��;��� �)"򱌬���<��?õ�
{�
���۞a�����T�P4T.�V��J��o�9�loW��U
f�̹����AEvo
X�tC�ᄈbfs^��L=gЊ:ٮ����D9�,��?	�>��={p����_3��5ļ���(�2*>CVI`�.ar��g�D�ߔ�E4�Y�0t��m���'j2�+�f䓕�<�u2 ��Sb� �a �XAPrP�j����WW����Z[�N�[.Λ����t%��ɽ�	����2���8�$L]���s���˓*Ċl���j�D� ca+"�+n�������'����:���}a������rob	;G�Ao��̎*�ƚ��Yr��xt8����.�ɔ���+��"�.������9G�}-˸���3�P�|<`D,!��],=522+����|DV��>`�o�uÜ�X�13�m��i�"}�)�����h/=u�>�U�n��s��Q�'\��&3x3�KZ՜�;�t3T�+��r�,�z�`�<�~��,Q(�6�)���a.m���?���OX�T̺�.�Kr�2��Џ
�k�C���5�	3�^�˨K��#�}��u[5��~�	��z����)ȼ���B֧qC4�\��Xb�aý�;���j�+����z)�z�)���"sA
���W����:�V�c����!
c����Q���d[�Bͱ�FQ�1�6J!�#υ��֥����F�x��X�H�	��IC$��G��߻��f�f�u]�Yz 2�|̬�#�(�H��٧��n�[1�6����Uߙ�%��]��/��qїb�8�����c�+V'{��:�&b�<d�b�r��{���I�>�B�����͞������$T9��y@\G&b��u�r��lo�����#֜�E�/�T�̀���=�ǔ`����W�;T�EZ�R��+��];w�˟�b�d�Xߑ*�Ö�J�e�\���
$�u�#P�ߤ� z�[�.�2��{tg�(+�*ㅦ�r�Yũ���	B�8�m�!A4�9�G�	|t�7`4$��y]���!ǥ"��Yt�h[��
J}�<�5W��Q��C�@a��a��ZkA;G����`����1\���ۦ����fN|
�Q��ʞcuAk:�
�eH�fw�D�#��x�C}�!�M.��a��xBN��r�[1$�����v�L�D�Kky�����e�?��.nƺ}a�
�������R�c*���7V|�~#��M�k�����X�����V�Tκ�����sŌuuX؛UY41���[㘾��!w��5��Z�D��/�#x�OC]7�^H����mh$�6f�iP�rOܜ�
QP��Ra��~��_�^���H�7ĕ�2g%r��<�ZC�I��,���K��꣟	f�7=Y�#�J"����8G264Mdq�XEXU;��4p���F��tմ= ��(]|UCU�j
%?�6��Z�,���j�t��UF��9A�y�״�qu-�VJӞX4��l�d��t���g���G�|��}?�?�x���Z1�a���q>�#��
e_��Y��qO��/����eG���~k��+y�y~�ɇ�mukڔM,O[�=�Z��ѻ���8�ק��/�g����Z�����f�k��#A��66����i�����
���ҷ�8��uK�k�L���㟯o��ꔭp�p�O��K���{R�zJ�����C�E�xÓ�ϠZDu���N���ϯ>.���m1���-4����9����z4_3*b��v���L�U2��mOӊG��v�\֤1z)�8ze��s���9`��k��U��u�}8嗢|�M�������N��z#��hW�=6�f���_H�}_8�N��xJ��a��4��g�'ŷ}a3�}Ys�:�S�F��-�/�]f��M5���ú��}�|y���N�4�XF^���&���pھ�z�ji1�X,�a5}����Μ$�P�1}��!ӥ;#��/t|x���𶭯ߕ�$r��ǧ�*������t�J%�v���t�)��!]=����{.>sIpvC,=4N��v��=}yC~)����z4��x���+����t��kGz�� �G�����D��}Syr��P�l�i��[W�7l���&�"��W��;�z��^�㸟�ﺞk��WQ������>�o����=�a���t�7h�ۀ$����;nJQ#���-�tM%�M�؉61IIF�ɘi���B��_�l�^�M��T@�$��/�t:����ܶ\��3������w/�������{�'�A���0t�~؏������������;�VO�6���{�C*��!�J�[>��`=� ��ّ|��ϛ��82X��)��te�XY�$���
���3x�J��X��>��#κdse�e2!cZ0>�SM�֟Y�ۏ���*��"�@ޏ�3���Ќ�vT�*�`ʐ��W�� {����_����o	�[�SK�H�>�-ww��{=�@{��`=� dӛ=+�,��A�>���K�t�*�]V���w���&"jS�R����]�Ck� ��-�]������Dn1�3�Q�,�ZDL��V��S4�t{pe� ��X<�=֯@Q=�Jq�U*A �i�z�L����4�#x����7�F���R�&b�@k�<c��G3�S��e�!vI,��+c��p�(�%((R3ܬ;�F��W�}����V�?�0�D�g� �����r,�Lk�E��P�
JyӀ�{-�u ��)lʸǕ�7u�{~�x�
еJ�f��>����*Z�'��D�Wf��ջ�M�Fe�@��x���r�]��{_��Mg9��Nj����E̸6j�&�Ma,]׏�wby*8+��P�����+��>�9�J.�,��<�K�8��³����}E�e�Gk���{t�
�G���d�ؒ�Kҿ�#�A:De��ƪ�s�S�2	�`�ws�8$��=iSLoC%�8z�3�z��:�0� �'�0ޭx_�.M��,t��a'�/j�in ۉ1��ڙ`�h'��o~���OkW--Dc��V���+�o�s��صE��܃���D �z��W��j��k�ei�^\�>�D>FP2i��ߴH�T4���af�Ch�bo�,��{5��ߞR��Qyx`�߀ڋ2�k��01���o���z�oO!�+��X��]����$�)���״wx6��(���Y�JtcE]"<)0�$�N�Y#&ŕǥ%F�ˎ��g�ش�������d&V���I~)=)�cO:>�xu[�X�~0����� �.^$�d$���A����8
�/�T��C����F�$�$&6�,IQ��r���6l�֥&���u.��'fN������[�f~�"�P0QDT+:���������'|p�3x\���5#^^���׻��#.�Q\��7�0�\¥��8VL�l�ʕ�d͹�;��,.F����C�� H��Uw<�B)��(��d���grÄVN"Ԥ[~��Y�Z��i^UQ�W���{w�qZd��how�}�])٤4� n��?T�#���h���f~�-R�vL���3�mA
m��t����N#8,�;őz���Z�WCN�LN9*�<���0�{�8V�t@1�p����GQ�@Vq4��Gd:�i�����r.�l9�5��M��IV	m���^8��{ ���PƁ��&��8���}���o�*kˠ�t
P�G�̠���܃���ӹ�羯d�z����M� W�)y��Ԉ�(�wY�p�#�L�i!6k+t#H�~�����t�Y��eW��:�ȹ��[��5Gp�O��W�p� %�l��I�X|����� �(Ɖ[�F��!E�_F�X�t\�ۆ;IF�FU�6�#�U-Wv0l���8���֣�I�	[62�S�V��w��n{e�nP��������$��
��0��Z{��n�M=9D�Hٮ0̅w��<c+T���h��
3�.iY�Q[.��}�޵)4~�	��suw�������c��)�w$��
��@��E&1o�v�k�op�lv5��nv�g�u-�l��(kD�D����;�t��A�]�t����y-n���l1b�<uخ�l]1�������5
�V�k�Y#��;��X�E���_�ex��P�����Gq�����a<[��Uh��&��cL��i�Nˢ�=����C*RZv�Nyi�8;��_Wخ�I�)�c���a"����|%�d�yӔ�M��Y0���*�X��{V���=z77tsW�U��	I����8��-o%ֽs�S8w�^8c�/]�wN+7�}�㶜���/v�`��%��x&��߯l:u�v��t�Wr���;uw!Ǒ�N�r�&��%{���ۏ)Fp�}K�:h�^w���t���
�rJYw�t͖.�eHB��h��<�����g�o��8��-�14ʏ.�)f��uY�>�G^vw(i�bOq$VƆap�)؉�79�$��%>|9�H�*��>�)w*w6�C�{p���e�x���_,��9�T�nۜ���;>7�����˖-۶�߷|A;�k�J!�R�oc}t[���]'�=����i͆~~��e�2!��:�PdE;x����D�ّ$$�F���{?��9�=��g������^��ݺ�W�u;߿�}ws�6�O��;�Uz��n;F�wn2���j����6Te�����49���Vۈ���F����<'`�m]����8Vt�������*v�g�8�|�2�7u�{���9�q$Np��{�{�>���8�^ƧbŚ���r7w\�Ȩ����:����-L<�	�ʽ�1\�u�`�C
{#X-3В���sUbhfY�=5zmU5A�� �)طt�)�4�B2���#��9۪�����&:Q�yu��#,1&���0��c��{�*{t����6�c͚4ʀwt���q���O�<.n��Z�h�m���/�M��v�fH�྽�1�L���e��x���B��Q��1�s=y�KVDw�0�Yػ2y3=<O75P�Nv�v�؝�n/`���Y'0���8ه�ˡ����^G'�
p�M��+-򡆺�'4LVZ�U7l�|��z�Vd�fD)�Fo]vYbg���bb�v6�����o/�(���(u�4���xȗP]D*�3Y�n���\Eu�|zZ]��W9���'%W^l�����<�ګ���
uys
�=̾B//4��5l�2�g"a�l�����Tb'���jsR�Юӛ�b{�� �9��y����.����e��!8mX��g;��yn7T��aX�J��TR�]dkӻ�K}�&����7�QX�%���&���^Wui{
�v%o4H�Û�]Z���fj�Y=�fF$��F�#\����s��T)��Q1����;f�u���n�K�֦�+���d�S�^�XX8�Ӂ}ss�.�"c����3�^�02�dQܡӸ#����3��T���d�yyP)T�fc��a)�6�"��;��]�ꝵ�5F�����9�����鮢�{>�3赳�}~�+ܫt���1��m���7��] �hY*�WMegLk���6��"2���R;//�-ٹ���̍�
��T9�W�I�3U����M�=�Y13amj�A�!�(����N�ڥQ<�X��[e��P�5^a��̈́6D��F�ΩFS�
�`M,���MljS�٭6��u��4J�:{^(y#�]�����LK.H���wx�͜f�'���{5O7��:�o�D힡N��&�m�{R�P��)���,鮭�uT�T��=zfjxR�w�n����Dd��Ӽ�K�!]l sh��9��5J�U�pk$�y���j���z,�Q���0�tv�=�%�r�C���*��.�s��<��� @p��x�W��nT	�U�E�Śt���b�"as�x�u����qM����ǅ��Ҹ�áaT�˱b4�����q�P�p{؃F�A���ٛ�nq�
�y\J�n������o�]�.7q��&�D>�s��z�䝫��6�ɉ�ȼ�U'��w�#,\�jI��d���yZ��O�%����L#�E=�"G�ʇ`Ҙ������7��)�F[EP�n�P��y�f ����I$m�����X�*!����Z�xb6\F	������Wu.�d�h��49��-r�6��7����2#_J�w�Y؝���%M�.�)r��*#�\wS+�4�*d�ͺ�{3��5#�N��ʉSmCɌ�6�^�Z�v�)B5'�b���w�ꋺ'Vs�u���!��n#Yڗ�Cov6��H�թjwN���7�-���tַ��BzPP����WXw�3֋��r�UuӲ����UͱoMla�+5�1G�║�U��eD޹b��!�:MZ�*8�.4�q�v��ޚ���i��OHfm����T.."k�B)��Į���t�]�/w��,�93�z��E�s}�Q�|�lS�A�L�S&뢱����j'�w�IX�=["�c�����S��J�N�X��o�s��}�b9f��Yy�� �]M+M�i꫇���s�md�ڟM���;A�4�f_��Y�͉J��c���a��������le��!��#��J��]�v�`��7�5v�0:�v�H�q���oL��7�3�Gf���A���6y
�I]�=%m^�� �u��w�ͥ���/�!�B��W99y=���M��:/dF��;4 �;���N��'1�$t�Ij7�����j @��N�iP�Y�]��.LU:�uh��bJ�鮬��ﳸ�)ٝ�ͺ��"H�Y�ɩ�]'Jcsye��q:)��P{���ҹ���R�\k��yԫj�<��F�a�˝WJ78���#DY1�p�θ��&�⺚���]6��e%���ܭ�-�tc�I�AB�<Ӫ���/��XE�A�9'xp��!I��d��k\�i_q�u=S�P�n�ʬ}6.�;:��� ��rC�������u]J�ݹ��B�B{6��rf�s��3-e�ǋ{�rU�ĭ�M�Ƞ{��1�y[�����!��$$���P�0�^�����Tge+���z�b�U�U1u3Ɓ���%��e]�*����^uu��Jp�$���׻t�o�%��`r���L��E]��]�y}tl�y�f�a��"Pٛ���Vu�t2T��%����QU�5j�o0u_�u�7��������1bqL��:#�d=��#�t�7��h�/6֌�{L�5j��n����w��"�rwD��+��J�Č�'6�n\NTN8�椌��=J��1�i�57w�.y�����s$�p��jc2宮[�3�;�����K�!I���[1�c��s;{/*'`ޗ/j����{�0�˹�ꁰݸ�Kh�u�D1K�w:T*�%�L{S��2�=/���G�ٝ8fh��H�\��q�A����%��2�$��%�cB4�����������uR�G+�+(M]T
�^c2��!�A�F��1�)���c*J�6��b\��7:/3f*p�\o%�Uֈ��n��v;k�a�V���@1���tf2�Mu���s�b΍����b������[7*��<Bt���z��Z�G�5Lv���Vw<ܙ�;'jl�}Bk�x�����X�8�	Xu��{�Z&�J�<���g��P�>8�غ�%lQ�۾��h���E�[�������R�2�ф����4��^:�NAtk0\��8I;3&�auY\'�w�c:����(ԣt����]�0ؓ�;:r1��ks�l��*�����ȅwyk�vfz�f�@�ى�5%.F2"�Z��hJL���}5W���Y&���78:�;��b0��Xv�+��bWe˱f�"�^Mr�N)�ʊ�3�Uɚ�����wd������0NI�ő�^l��/�d&-��������k�
s��ع���;ś05;�=�tOn�U��u�fG�:B:f�㔇�Ft�g\�s�Lj��:�����'���;�C<vhP�0fl���"8lGK�ʙ�NU5��]`<ɨ�s"�V*�R����N�죬��w�wvv�v����e�1v[|vw�d8�]���:&{+�H�Л`��f�ޘ�Uĳ�7�5]���kgc* A\�юt��Ɉ��Rv�eQ�vv���sS��l%�ӵ}s��qviI�RgD�0���u�7��g:iǓ�7@�"��o��ݫ1�q�݋O'jrheOy�a⬭��������Q�".��ڹ5'fq^�)��B˖fg6c��r�2�Kn��ѧ�q�.'#���ۻ��`�B��uy��(ͱ�D�[�DJ}���K�j�f^>ӱ�R3��kj�݇F�OFwT��'�o�v�X��.�:�������+I羡�Ϧ}N�>�F༝ݬ��+k�|Y�5��`��X�b���nLN�D ��M:{�՘��>�͉���j���[����/��������W�s�v.���9O*���a�=a;3�el�oUtb��S@I`�殃ʹ{�OBK���U�%�Vn3f��*�q4�(�Y�92��lm���[W{.g/Z�UQy��WOn�n�l�7���j�W����u���ۚd�./n�=.�&�����ƈ�u����'C��JQ��8���%^C�}1ѽj����Ӥ�7S�^U��p�T.&*�.n:�;�=�·*�f!�4��A\���ˍj6j�n\Uⱪ����Q�����7_X����.}���=o��uX�3X�"J����wb+��\�Q����C!ź�k,ۍ[��׾�׹�nG}�ݎ��7���k�4Ι��H�M���e���O����'e�u��MO:ۼP'��g�6�1f�hW֝�UWo�Fv,�EF�:�,�"�w+���U���9sę��R���7Y9.�I�K&����^Ҟ�X��==0�y�Qrk�l+���z���w�Z1�օW�{�EJ~wpo���-���j�	�{{re�ޗ�Bn��&�bc�{���ی�4[ĦYt��:x�P�Z,ՊIJ�e��N�u$��A�4�׷ѻ�����g�a�.(^Y��ۈ�����`0bz�(�茌�f�b{y2�d�:��ʞ�n]E�DQ��Cr�W]V���1̧/�����}B��5׼��#'n��;Gj�6��e����&��Ks:��p�݄X�̑��g#Q�odapәT���v�;\ў�`_pA˛#67�-�=��x[�/���2{/5�#_��ݘgj�V''j�����v�
k%
֢MU����1���.�'/�9�PvU��j彻��qv�<q̝K�uѹ9�����g�)�nv��p�_9ײ��78�ܲ#��D��Ԫ������U��;d]S566�=Ev9od��P.�W#z�ջ��r��ɛ��Sw=m�J���l��
�+p��<R>Pb��+&.��ݥ��S�s7��vbe�.�V�5�3\V�`�5�=R�:^��_B�Eֵ�ڻ��؞V"E�wI�[���:���e7�j{��=W�tvu���xomU���*_�nԝ
j����z"]�cۍ3�RT��P
��tI��y�N��y�Qy��̃&�U왵=/z�b%6��f���P�;�������1��c�3�c�*�T���Øӱ{�+�ȉ���xw�9b��*q�7sr�!eԽ�0�+�8�b�R��ܵ���]2cɎ�OѼ3#8���ὅ=�����v��N��*cg(��������,M�J�Zu�NU����T�����c��Bf��":.K����'�7
¢�$�*�r��:�S8���n/4oc2�+��Bu9T����j��k[�裗N/&¸�=�s{�|n�v���۵�h�MJ�C��ν�Rg�#m�ܼ�*�Q�5r�7�Pz��̧�����<��^Y��sY��B�*�f�WBu���f�b����TH蘞˪Ӛ��CɅYԫ�SlD�����5Vl�n����w���};��8]�Tn��oy*��f(�eZ>dݗְn)�1wq3��uW.%^�o��(Yqu��v�ѡ���O]2�f]d����q*�L(�ԧ0��6t�ܼ7����ɸTr##N}6A�٨�7�edR��[P�No#����ш񾈩�Y#:�d��^�q�F�Љ�Y7ٮ2|����TT�����+L�{u�[��uƚѲ�mT6`��v؋��]��2�r�z�/F�c���1=1;!�4F}��N����BA����צ��fk����\
��諆7\�#tmܨpjsd���=8�*���'��}8^���2V��l�^A{.w/�(J�'6�ck��B:A���K\ɪy��{!N�Tv�:+}������G�=��Q�OUF�f�Kݸ>����~���:�@���5u������5:d�������O��UZz #kT�n��9X�͍ۤUd�ɧ�z:7�]쎏k7���o���=Π�-����;3xE�gN�v�͞�7F.uԺ��:rv�:碞]��"5�ýz����:�R�sg#�u^U�.I��ULT`Χ{o���=����;���D\�����&�e��y!`D	�ژ���]-T�Z{2-���H�g��S�K���6�v�ɪ�;Ff��y(_z��6_l�-nv��,h]�:N���b����s�Ĵ�fB����F񬋻�}���h���,��Ǳ�n�8u�J�jh^�S�p䛕�w�*��X�՘��^Z��YQ!S�õ1�c��ښ���c"�LP��GwsqVM��˨�z�ԭ�����suЕ;��L+ڈ�{�Wp�Y.���Z�6b�X��t�6�_d�Xqt�S9�6��8�'���F(��اL����Z.s��Χ��%wYR�b�m̙�c���%T��|2u��w���t+t%�e����f,��sw���/I5�'v]<�Yh.��iءTˬQ}��{kk��ӡ�8�{�%�D^rf�a���3���p���.��E<,v���z{�9*}����%,=��
��;ڮ.�ʌ��ݼ�+X��Q�&�D�W3��8tm(BWr�c!��\�mtNk�T'�v-���6�c�5��p�r.��ێ�Dmn]�b�+�bH���a���y4�C��ݑmO���o��P��鳹q�&�Y�^���wӫ'����of��oT`���A�5SSjN�=��V���3Qˑ#:��*\-ޘ�����#,̅�yW���_�pS&����j�gC���2c�$D��Ya�Fe�!�6j�m�WB���P����
&�dOF1��-��;+�����f/d��Ebˣj߲��Y�O��W���T��ȩsoNwF�&���Qv������t�j��3�Z�6l��3�帖�E)�s�p���͑��h��:v�&xwa��=�.�n>�8�n��j����n�u������p��tM�`ŌX�6wc3j���sl�/u���{���S��:+���1F�)Sf&��E��0A|����쥑q�^�u��L�T��=�y��My{�0����&���"n�ȧ&�R�R�$`�ɉf���^䌉\�9��s�{�,�[R2(�A��L��Q�w��E+��ԩ���MW�`'v�r�=���a����˷�X�$|�F�8y�x�Wה�Ԇ��i��u�/�!�+pU�q�r���gu^+T�j�'pE�����ɞ\I���wD����rצ��z*��42��������O\���/�͠v�*:1�F��>ě�M����s}�z�:&zjw��l=�^��g0�S֐����.�^��+D��ڽ0���f���-�P��Ӛܝ����0�ˎΉ9���"#�����PoU��^1v՘�Z�S8As�fg�D�s10�dZ��S+�W�&��Pɴq��C&"�kѯ&��p�P���81�nV��qM���@��2����JW<�"�7C��%��=�GwN;�p�φa��e*�=���u)q��&j�s���:̙�%�n�l����s m<�֡�}�Q�Q+��58�Kw�U
(K@�Q�[s>�O�9W-�h��ѧs.o�T��3�j�v�s�EAimOdf�c��ͳ�+\oR��u����D�i�o�_�]�X�[�r�}�u<�U�g�(d�Y�/(�X���3��Ճ���˵�f��mV�v�y%OWCp܌�Z��n�spG�s2�zjOq(���^�[Uw�&��0�[��V��-X�uEn��Kkk����Zx�!�X�<;q�Y����E�>��g8F�w7���3�b�9�ۏ"z&���bb�c��)A����Ɲ$�9�J�]q7ѹL�Z=��q��퉨�q}0�]�K�����Mw�Vz�v����[��Ĕ`�>�$n�W���N,مa])�!YĨ�$�k�_�2�	���w��s;u4����#`�$�c��ñ��u;Y��CzU�ky�rc�~�y
(��L_��n�������3r}αO�˻���c}�&&�n����}�M
��ޑs�������V��hB��Cin�^H�&�.�,�L���Xo����Lw^�$od4���f?6%�[&�x��˃���le��L�8+!��ݍ�G�j`ELfq���������t�s�ge+E�5��c�&h17�3:UU�{zzt�.��en8sJ�=��n0���j4����g�w�q�w�15R)��R��c#��xU�!�`��אM�VU�J�#�T����j��T��L^�>]lΈ�ׄv�Q4�pr25���X����ݞ";�5DvFI����{��Z���k�EŒ��e�AZ��ʘ���h㸊��l�|�]2�"-�9���p�=���{*��MY7�7{ip%-��p����.S�s=K"���/�1��g+4�{$N����M�0��^OM�ݥ�k%Ց�*&�F�!O\�EONZ��;��ud����d��+��Zضj��S��nzD�(I���v�X�s'�o2�2.N�:fح��	�;lf��Η�/����D+���*�Yk%�]�ѕj��gI��y�ػ}���׮B��*+U-�LH��n��sy� �����.����̓}���[0�f�D�{���L�H��O�3Qv�v�0c."&'ۧA��m:걙�\�+d:�xL^g[�ͮFIy�;�.�^����8�٘K]U�
�&7XQ�,I5��kɓ�.V�@�J��(��3���$`��Z(Mf��!����7�۵Mu3{��l��ȲFd�U���[�4M��I�ʂe�b������k.����r�V��Gd�єh�4��M��{���tGq)!�'�D�b�'X/8V]�5���q��t�M�Q�=]&.&����:��X��4��s�q�eu:�r$��e�14V�R�{�q�T�v�M\Խ�[[�E��rflp�̠'c��Q���黑�{���������^xagD��m�͜vnd�F�[w\��rvĻ�n��
�Vl�L`��1\T�V�[{1�㵼ef���Gd�M�;�g[�wy�o����D(�&wg��FZy�;�1ܣǺ�0r����{�-Z�c���J��tFM홻��}p$2�ٹ�11��EO�\��|'�gu֞���F�O�b8X��ts�d��6P�Jᛃ]���&�Fpw.�3+b�=u�ƫ�tX�f�U��<6c,�:]���V�;d^ܭ�����l�)�m]���#0��$�uʊP]q��0v�X6�s�ت��"��/���׮��ս2��U�ZmW-W�x��۶\yskD깍�qwӸ��EqQ���/%���A�B��o�j�/E#�����w��'o&���F�%汶���u�OGK;\��M궮3���s��&9��*�ij���H��X%��NVn2����>�����,�l��;��1}`͚jq��`_]_WEӢ}���7�G�X-��"b�Ӹ�j��gY~�噜{v_���}p���N��諦b$��nrD�*{�V��nlk0EI���e\��"ܦĪ�==�{\�Rng�p$��X�[uO��+w�F������s+����3�|{0�f�ٺ�yI��8�
!Z�s�]ٱ����!j|;D��ƪ���nzk4���������P0�Y��!�G�NK��p�}���X�ۢ
t�&�'�!K�"I=7�� �f����J�Q�a\L�0���eZ���*I�PLM�8�a�y���Ø0Ϙ�0z�M���z�nddS8���v{�(V�.�J��v��]��0����I�e���z&s4��qw��GTUm>���x{�ěXT��j��+�^���O-�t��2c�K�1�+Q]c�E"+�Z����a��j��]<�2�m�US3qBI1ӻY����Z���WJ��5��&v_fA��2�+k�2^܈�t�������_M"VB�y�t���	��'دJ��o25����ׯQ��0��3�r�l�8�B�}�Dg�!)���sP�UL��]�f-bx�GOE��L�طLeԙ�|6��r���7ȫ�MN�F�@������-y9̷�k]w�n,=؄c0vֺ�lB��7ݒyqɂc.�E�j��yD�C�#����59]�1�f�M��vVT_Y�M%�a5,WTThLHЅ8����b(�U��ON��ٖ�p��qk����D*�]�71���;;$���7r��7G)`')^�Y�cd�SO;\���v�H�¤c�g�F;fnn�i��\W1vቶ�^'Dr{l��C�ԑqU�;�e$G[��^ѡ�6�3�S4L��vC�[���{�07a���AY&��ُy=5�SAMh�h�m�{��ތ�43z�
9<t��GMˢ�Ȓ�ۭsB���c;k�b/ngT�^�F���jz��9&�1�42xX��@��9MguѲv����,��ݹ�s�����j�7���U��,WN9��b;n���=��r�T�T]c��
j�/��ܽ��/�@�W�4]y%h�:��Q5���V��p��(�d4(j�`u��h��Ү��5}5��Ϻ����9e�$�b�t��U`�5���jܽ�
/ܡ�.F��:��II�7����{,��8��6�Ԯo�8�%�!K�C]�Ģƌ��rT�cf"�$rq��5EE=���3��H��!lL.�,{*��HR�PT��K�ELYq惙���V$F�.m�T,�Ѫ�S[X���#mi6�q�ٱ�K.��9٤���Jl]��쨭���6��i�-v]�����MCr:iwsk�č�&#bB�v�˹��0�.�İ]��4m].\�����آ��u��EF���*�뛥	$rܷ�F�F��K"�v�)��\�.��ˠ\��H�D��ذ!�"�7�ҝ�ӶI.h�!su(�gu�Cd.v'.Eҹ"�ݚi��j.\wQʃL��{m��U~��m5ȴ�SNk��}ü�I۷����m=�/�x._��\M��?}���e�w�� &�G������p�̗�;���Fd=ړ���{|�'[�@v��]Z���7/g��>[�W���7�f�ȳ
r29����d��V�'�����[���!Q�m�!3���L[QoK��8�A�'�"*��-�o�^�+	�c°�5��0�����]7`l�5�Ud�TJ�X�p`���9��a�@����l��
�~^�h�F ���sCb\>�����Uz�X�����i@-�V�wv�!��2�N�T=GB�03�����G��)���O�N��Q��h
��'�ЂK�%鵏�^��B7i�
՘kT c��|��kTT�gn+/&�J�f^�pߦ��0=��k�\*:�9��1�Q�k���E��, g�§��a~��!��Ê�b��![P���5��:C6�O\.-�zr�n�¦vI��(n�ǌC�Na�K��ѧ�����v"=�T��x�Fԥ�Ґ'��,b6#��%�T��t�%�|.ύ�hw�ԉ�r�2��fE��J_�?cl!S��|���a1s�P�xXV��t��!z��Z�0k%*L͡���؜�O�W�,��r4���6���1���(�v.�pP��]Ȅ*��>N�ev�z�C�R��}'jVM����2��j�W�>WI��v��=}s��8k�)罭�wp����z����-��Xt��=q]Ab��:7m�A[v9%{�!��!u�|���Ю�'s+��%��O*�A��e��zH=�Z�)���/[ss�6x�7A�Z֊F��?&鷮�ѯ�"�ε�Qh>��i��[��<��X��^�ס9kuE�f�2� �&*���!�z�Q���%⅋08T�jW�;q��dl}x�<�:��� [Y͔�*��WY�����g*���^�ؗL7pZv��ñ1څ�Yc2랝5�V9�5)dϩ�!�UIW1wN|�s��.˓3$���s�\/���˴���dr�7Ӗ7?ٟ^���d�O���,���N�x�*|/�żG�dhu+ v����B�8�mC#,/�q�M۷Ql�p=_�5��H���ٽ,�\]��F������M�l7a��[���"S��Op�ϭR��Zn�J�饕Ѿ��[/ �.Ϸ��	w�p�a��a������_�-P���?��EK����ٖ��;K�
xΝ?�E�Ƒ��亥���۪���;g������Hc��>T�����dk�g�uLL���J��q-1������lq�����I�a^���-�� �{��w�f.I�4�lV`<����QCʺ���&V�r�x�ј�Չ�D0t��=^ b���͊�)����f�*��u��X�U���6����1�]����J%�~��Lr��3��O�N�T��V���"��v��������Dj�lUr�p���5�1$�g��-4첆����+9c2�z�`Da��I��M���9�oE�a:ܼ.�k;����c�J�_J�LnW����V�J���E˚._�{�)��B �� ��_~s��i
��Ɏ����hO���`�Q��H�P���9���u�
C�fyj�Y"��1�§脶��cy���;tߌ���HK'�|�D�N������RP����p�%¦,���`�d����T*vz�����=�qB�C`�[��'�2)��1��IIzr�ԋI�ci�c�û��x�.�����,q{i�:��"]m��}5 ����� =��0��nK��w�� �a��n���w/�}�8�mU�խ�k�o��퓼�[�!ͤ،�F#���}B��1l���u�+��{��ۇ(�j�x*[�Vr�Rye<�3�����ψv�KDa�4�x?J�aͮ�Ǌ���ÚfE�9m�<�9O	.s�Q:��ȵӎ�����j?�<p���
Qό�H�t�����?r�󽣄�\��^���+h6�L�w��q,�U@O>s���:�A�9�{i6�k'L��UC�Y�t�C��S�9�k�#S
�1m]��ʸ9[$�_,�<i����U��R�pW���|���G7�j)����+���q��l�]k�8@a�>\���b��^z�ME0^j���!�0�8豋k�=��X����<����y7���q�x��k�7E4�.K��vC��`��tv�ʸ`�Ƽ�o���Gf�%�B1!πȄ�09���������{O���F��}O��}������A�w/Q�:N��>Fh!� �
6�(	��6.��Dv���>�����=���_s�a{~W�~��I���K��)�-��#�����>H>�_���)��/�~��1�T&9ٵ��_�C�[%/���Q�}�ICT�o�*���l-|�Aۈ=��bW>��|�+��!�*|w��W�]����D�f���M�>Q���k0��r���{�;V�o��}����d =�]4��������I2A�ѧ�t^l�iiHD���/ɅP�w�  �Z����B]�}	�*���.�g�P��t<��\#Hx~��o$'� ��"$ᴲ�Ä�����Q7��V� 3�h���v}h���-��C�r&|˛G�&ގ#�{�5�j��!;�n��_���7�L_Σ�3�ei���s�1�/���ꃤP�qM���戚#�}`_n�ø��O8 Ĕ��ь����*-�,Z�N�]E�C	Ҡ��i/0z��7д��Tn�^]^Vz7��J2��So�Pۢ���3�Ӯ��c�*l}l�(�S��b�\*�aV32�<�v����p�(33%&29
���]��=<�C�"|�f�P�TD����#ڻx6��d�.���[�3�����ghpx8aLŇ�'!*�����R��]�r�5���i9J/a&1��ԃ�y��dЭ&'�B�;Tt@;5�i�����^rB����C���n�*kŹ/Y�Y�OĞ��)�hL��-v��ڏQ1HQ��e�d�_���t��[V���k��~�s\�Fs�d�@a�%�-3f7FBz�AĠ&�i��y��8��(UJ�f,*J�М����V����x�=�rl"��u�bǬ�P�&S��߃�j���_�|�{s���x�I�+��H�SOM�E�b�>ĤТ�R���}�M$�Nb��_H�}��Xs:fKu7N4 IcőЊ�2'�M�_(��� �G��YҎ�A��'q	�V�X+d�s˾DS���qW��M���GעEI-��ֽ����XW������::鸵�xv.��M/"ev4��s�
p�3��<��@�2/{��eiܫ�*8���t�C�.=�9|#�<Dj�X���F���=��_�eI.�l� Rn��v^��*�	ϢjNJ$�)V�Ӛ�&�Ig]�����cϢ{Z�`����Q���[{�Lt�b���,��=��a7�W=I�=$��`�bkru��k���e�#��l��!P��=)_/�i�TB�[����OlDG��4�B��|�Ġ������P+K/�\��ceN&��-�{Ba{��k�y\3�͜��C�D��%�M��1�sn�M7�b�Pw��
���v�
���bY�'ƪu��&����&IJ\0��ZŞL��Z���ӻ�LmwF���l��W7�w1	�`jMK�d�Mdv:� ��^qTGp�r\,x�L���Q^W<,X��I��r?	�;4��Ue��x=[\M	[�ʼ;v����M��@�8n�[~�^�����G��`�Hy���dR�jk�k���գM�SP/~�y�V�u����+��N(S��kT�`�QU�S���;��lz}�[�=�OF G�j��Az]�c�s����盥�n9V[q9f9�q%��On{�{u��v���|�c�x���8��+��t�Ϫ�R<�����>�C�x�K�	2doe��zᆕ��8���y�|ʴ���ځ�D��H�K��t����T�{7����|'��҂G2�9�S�FK�=�:b��������+źc[��g�	�o�q�)�ǐý"�{�<���]vО8%�f��cN�ܟ�^xOQ�����s���,�I��������{=��|����_�m@�~���?y�g��ݣ�	����y�"#��$�&	�L��D^�r�mm&��$��	Y/��/���-7M3����Tf�$��i�YBj1�Zg\��,!$jB�Ͷv�4{����M'�ۼ�D�r�����v{^��N������I7���Z^kUAL����Al�o����he{�Լuz9�����7�g�Z�a��,���dsHD��R`��~vˢ���*�}l@���g.3�L���MK���l��2P��Z��О�w0��5}t��M�
n�\�{�A���n;�7XZ[�s�g}wP���䪍�U�oj�^K6܍�ݚW+k
�	=h�8g�b���ޣrK`�nU��q���{n��&�)��ϿZ'yET �D��%mS�U��X!1Sڟi��?a�7�n���߿��~3�k����<W��z>Oa��?���vߠ���ݨ*m}��_�ykZ��N���E���W	�p�.)��=�n���ٷU���E��/�ǒ��y$6_�9�+^�9��囆H �k��\�C��9�Dh�Qᯮo}WIZpp��⋞X9���e�HA5d�V�Fy���8U)l�Z��N���b􊹪ֶ�2s�g�x��L��0�q6~W�f��d�k��X��b2�#>�v���}��q���p�Y`�psʆ���k��d�ͳJ^�^����2���նDzf��''0����ܡ7���L\��+�9V��c�j�(��APaZ��2�UGIoD@��rY$$�����7y�<��Cu�}_��~�k��#�7^��v}�]�8����u����|���޻���O�7pB���A�D��� +jD`"�-��5R�U��[Sl�� 0@��� �y����w�����/��m���t��(h�z��+��WѰ���.�Vڈ�w뾨Γ�Y0��*��>�_������4��̪��LơG�n����9���>��w|[�i��@��I�����	�K3�D/��">�Y���J�~���Ó�䏪_q��;����SC���ף>_s���d#(���q�{��y?]q~н��V���}PUW�.b��g`.�C�
B �.�!"Z�v����-�������e�:���s�/�z�q��k��n�}�3�w_��>'E�>���w��W}��~G�?��AM�+�#G`���
U�"���m�r��_t��5���r7��_j�,ԑ��\)n����ApV����$�P���&�r=w%��Zܿ+_ga9�E�(�����j���Rw7��I����2�|�b7�^y2x��|긺c�B_.ǅ�c�R̂�"��93T��>����p�g/�����?���߳�>���~��9?+�:o?�����?��8����/o����S�[H
p�8����8��	�e���&뛾L�2��i��q��B�1ބ��R�uf����r�}����ּz�g]�n�Qj�z����DH@B�&0����*�߾���5�z~M���^���@��,�F?G�w�u,`|ߌ�sc>�|s(@=���a?$����ֿ#�k6�Ce��ݠ�.?ٿ�<���=��OZ^�e �Td��ty'o��͏��YE��XL#ݒl7�V�9�o��~A���>D��i���9>�O{�M�O���'���>ڈ��Ϭ�g�;a��L���Vm�-kf�Rg6CB�\P(i�Z�L�xO��4
I11:`��������lAKѡ��^
����
�Dxi&��EG�S"5���y�:h���c
6�@�~�4~b�-�XG�	�d�!yZ�X��>�n'>���܃lP8Yi2F�����]���I �{ebc��W��E���| �?���I~��`�_��5Y�g��� K-�I?�C��Z�Fɂ� �C�
���E|d(����B�l�z?�(զ���#���LP$��9,A)A!bJ?4���(A+�@��TO��A��O��d�Z�d���"���w��)���U	��\��U!�U7OS~�376D����j^�-|�����OJ��9y����'	�?�&d�@��Kr���A�h�6��Ca,��FTϋ¾1��H�<Q��n5��� ��T��pI0]���@��?���|��HDa�|U��LP��2��9�8�
��� @�����ۖ"^�UhkBo�������BJ$O��ϟ�?&���G��������#��v�4-!�Q�����D�3�TĢ	6��E��������^S�LJ+���T��"ɵ�0A�?S��h3��� ����TL6�����-U�D4��%����k�XW�Ԇ�U[Ô>s�m�%�Z�8�|3�&Lzy�ҥD�X��ؠI����mڹY
8 !�72�$gv�T�[��u|�
��Af[��.��t����g�����\C$2 ���qfS���5EFe�yc1�K�o��.(��K(��Z�V�GBE����Թ��- �X�3D��!�����*�9��C<��)C�R�i��5�\���$�m{9�$��(tZђ*�Wr���E��ht ���!�#`~2�I��}{�|�5��F��!鈑�+p;�	,+Iԧ����?�z�s�"`G��2�b�l2E�ف�+�V�1|�'6#$���ӆ,ZH�$�H4���r"+U��ኸO�,R"p��VC�д��ģR��e��S�=�迲��ꘟ��H�O���\B�c�}��=�LmiQ��Ċ��`��Iw���WB'��Q���G�$�$^���Q����==o��>a�ga���.���7���R'2�M��Õ�(����D���>����С&<>?���" �oFh�O��h%D�Zh���y �ԈB��b;GcTv%�(CK����K1�?	���d�Uơ
�u;#��zDe`��䀈�~�ʬJ�>Rm7���:<�����B�R �g��}��0�l��IkI�5�$��3���Ȧ�}l��r���~��}�>&�<�(��U��>����7��|5�`�'��!�4�?e��c: %X���s����MM�Z�ݏ���;P�����0Z��rk���#��g�Ht!JB�rW�
!ȀR	��
d�ϐ�B�H� ʏ?���;��0>�}H}�����?E��!�DzK�z$��~1�D�x�v�F�I�W��BM�����C�14jc5z�c��@��'�=ʊ֥?����(3,%�{��Ua����k�v.�����iR(d���2���v��.��F>ȏ�@MT���O{J%�|��2��]91'��!��߷����o�.a'�����|�ϙ���"a�*f����<����������Ѥr!�7o����Ur��(����3�<a~�e$!J�r잊S,���ቻ����1����Y%��7f�,y��.$o��8��d�vY$�?��u +@Щd-jbq5�) g �&c�$��\���>����#�'�S��!�:O������|@tu����6,~ďA��X�P�%�a*Z8�g��T'��s7���V0{�B:���Z�Iñ�TY.,'db�MV~%����~�{����y�ű���@�v�� �����F�!g��~��y�"3��������D�n0�(��@�<ߧn1����U��z$�E�&O�תNz�������wq�ڦ����%�ʔbA E�S.��[S\-�]0�Ͳ8^��% ���?4��&V��v���e�}�	}T }A��~{X���sC���MQ�i���PL"gtx�z��QQE�Z��lD������D��(*0F��ǣ�4y���C��H(�oW�ҡ�51�0+�RƠT�VL��#�3'���B&p2��pВS��$�0F�+<��k�*JRdF���a���T�խ���]Uypx�;"������u����2�m��l����E�=�A�����)!E(XK;r'��/�d盘��ȑ"g�Q��B�h�!HB�usW�ߡ����_|#�>�/	�8>�N�C.C���z�	�>X�^Y�[3�~�w^�^�����tI��2(��c?��0>FXﺣ�����J�! ���(�?� )io��1e|i䴭S?c��ۿ"��֏b$�q���- Bmמ.�!�P�������I����Q�Y����q�Zm�D+:�E�$��8�`T(����zQ��B]�H텀F%{a��=��w��>Yо#�eOz�'�G�5��>���E��WA����Y�I��bђ��I��
�+�������pS��r(�M��>H��߹ᩐ9�B��ሉnR��@�b�<����{5���K�ԇ�c��. ��2~�|����O8���/袛Q����r`��z>�+�)G�и���p�s��їZ�CE��kU\o
C( ��9�2����c�Zو��b�@��Pc
���u�Y�$b]�n��c\M�G�֦�5PI,5s����O��m�B�������T��z��f�����KLmF8:caG���28v?��>�O}A��P�>}�'<�3�a+�������6>^�O�Gʸ��M)��s���N	E[0�pG�j�厁Ĉ�!Y�Ed���bA,���N`�6��7�s[D��ჂȗQ�zΠ�c2+�ϱ ���ʩ!��>���������G�s䍡D2R&�@밥�8
��#�QC�'c<ci�@04��@5$:msh������u ��>T/��hM�𐯺I��|�v/�����c�GA�$���.P�5���S�f2s��P��-�(El��@%yc�#��?�|?_�AL���Xg��Y2���tI*&OCD�a�)`&����0�)��ԺH�l.�aAIh�Hid�>8c�3�/�� |qOvO�?MäAa�D�-�ʖ�Ԩ�-���@Ծ5,��i��E��CZ�7Yk�H38�Ld�%G=Q�MlubX�Uy�
�	QX�1s�Kʲx��I������?8��^��Q&�e�ЈV@-���ʾ�3K�q��심�|٭5�(�Ys3� ���X&�Q2&2"�h�T9i"+�f=���|4>|������i�_��	_{��;��+�޼>	 ���g�4P�@ �A�4/<���4Ǿ��z0���TA���A@E(��B�0��D�!P6aF�Vթ�H#��p�(B+L�*Ef	5	B	�B�H��:�սD"�D#�m�D��g��W��ѧE:�������j�^��K	�D��Z9�&����ȓmUQ�V^���A�B�b��3��>r�
(��	��_,��<�����b�Tcj]pk
�s5V�.�L\ĵD��$�ZP9*�#�U�Kp�*�0�@�X(�Q��`#vb`�H�U����>5�*Yf�a�y�]�4����n����&��=<C���X?[��H$H�I ����G��������
�h�Y ��-��Mb��&�D���3G�֐	�{�}�!��;��<����ݥo�D�M��(X�ޢ��;�C#B�q(�<�� ��dl�1�GFa�$H<��e(���M��|���u
I��"Q��pϛ$D��X�$�*���4o�I������^��H� �Rz�$�+Im�[X�#N��9�VTD�up�XH�
9$�6�VR$f�� ��ώ�������H���1�H> ���^Zf����"���
�����FA�����^f �%�Scq�g�Q�(�x MP�?"ǒA#"��ܹti5��W9��4� 162[IE���4a`B��"��zw�O���x��	��>���c���A'����		�_?�}�����I �=>I`6Ia���6��I%��\�Mh�rQ�F�����@�:� ���G�Fфt��LY�Ʌ�Y�fXFI�2�H�̗hav���.ɜiӳMI/3�Q*�(2�c9�ԁ1L+@�1	,ml���G;���;���H�h{���va$���#����!��Fl$:^��$(P�s(��1d���)<#Z�T��ܫ1�as�&b��.a���7堩 �$dX.l� [LU������W�$�+/IA%�������t�"K�Y�bY)')�%�kPɃ��ɳr�YbI�`JPcV��q�´@E�LMK0J���I�5sq�XH�(e1&am\)���22b~��a�/I�t$ �B��8�1O��#P��~~��� �$/-|���$�J�=�n�?�y��l���3�O�$k�H���Q�+�$�Ϋ$n��3Y����ӪΎ�0��#	t�!!���!C�.鉒hE���"�OB"&0�PA�I��O��3 @��!~��H_��e�{�h Bb�����;`��(0�v\�ʐ�ٶ(���	��M3�E�:!��2D?��'��G��6������(� �AΎ;GRa�]����Vϕ�FI"�����$�Q)zH�[4�,�V�G���Z,2@,�H$w�̀ekCf�����^I"���F�$�	�"@ed�� �v�Q@$&e�8��!�����ZNEҘIHI-��fl"t�D���(�L�� &��I��dYs�Ɵ�#��@#���y�:UR	b��2�o;�JS�T�%�\2[��,��Fs��I���T��j�'T������n� jY�AI���3�
	��4�9��X���P���H�I�븒��Z���JV�/�h�YN�q�ɝ��#��~}|�R�5����x@>~H^i"||X���'}_{��;L>Pq��>�������ſ����}� �A�`~�|.ސ�>SCA$�>�����H���_��H�(�Q����uω>$� �`�q�qΜ�b@����'�gn!���J	d�|%���G���=��w	�mPX�������	�M�e�� }��|�R#_�#�E�|(�0H�=�ܤ
X-"J���$\g��.�Q���W(�- H2}!4�%��L~_y����L����<Q�m`?�^!B�@$��� ��#�~�X?f�1e��0F~Ō�YT��d�����ǽA�?���Q%J�c��������:���?�I��_�������/��}Bd�����|H!e,�u��/��ׄ���=?��A?�� ���}6>$&A&S���U	BH,cE�&��߀�u������a�S�L�a��j2|D�	�h����6đ$}B���������_Z�b(q	�5H2�����@��R[���l�22%�)x���P<bJ�����yv��e4�I4�O��K��>��i&�v�_{��Z5�,��K���C��@C썊 ���3�,���K�����aZ��_��h+ꞡo¼�0��+�R B�L�K����*����K@G>���
D���g��o����Z�4�{�)A���`�%�@���d$-��~1A8��Q�&�b3�kJ�ZZw&IP�����ϨV4~G͉���"^����6�y("�
�$>L:��;>|߂u1���
E}��p�,�|���Ӗ}E�iE�J�tݛl;_�e���@�0�lȡVV�`�|^G�0,)/�!�H�C�Lb?���/bl��ƴ̶�3��� }P̴*�����~��O��߂ŁEO��� �A5P_���vY��%4�/��Z?�s#�/���|�
.G�~2�	4����}�5��m6���y!c>ДCH�Hh��
 }�����S����}G�[�����~#����v+���B"p@����{��?6��?/��$!��`j�Hƪ��ȣ�^[W�f�$�Ə�ooZC��'�|�(/�>j#}f�f3T���L��:��d\ZO����H�@��~�F�R��G���$���Hc�4��?~��:f�!���D�ۖ�h2���k�7'�C%!U��IϺc0���W���G�����0�#�kS��#慤Ym��^��<��R���o`8�-u��CaO�3k+�+'��n���L�&)s�����g|��Q	�ډ��\�D�TY��{���*�gHQvjQs�DH1,B��8:�?�����w�p>�<B� *�^*@,�H��� �$̶(#����Hۧ�]��F�L$~W�����������~�S�b��\�BR<��D�J��x#J���$k�s��;����k�O��$���[f9D4����h�$���Fh�*��K���s�%~oc�"�EY���E��4,�����!(Hr�Qt��C�|�s��E�݆���H�����^�& 0��jTM��^�Ѓ$#A|K�?��u48�㌣��^�>��8��
@M�BBP��%+�'$�o7�4���/Z3�� �������ߝ��}�$̫�!����畄O�?�h���;���>�C��Bs�򴏨����~������U�4�_�����
!���SQL��q$���|>��ѷs"`���L�?_�"������"�|�$v���Ѹ�=�L��]���?��ӄ��\͉��reV���c}���j=_����l{�*�}~���z\2K?��v|�� �(/@��3�(�_�a�(���K�o�O�����<�[�j�mZ��	Ż_g�Z�%��z�ʐ���B������?_�Q�*9��+���a����)��(�)��>X�3�@�lt�Pc��q;�B��e蒓Z?�YhzV+. 5��� �L��k1\���o��@"����4�^�ׇ"8�.�h�R�A��8�[��-uG��VDP���3��M),��\���X��7Dz%E�ev~�����6G���,6U$o�u���^D�3���Jq��2.xB�����
R�7���1�0L���Z��7L�.��$���1^C���� ��U��0ّ�S����[d~C���|����S�9�|�~�<^�")̪�����D.7\(Ny�ݍ���A	~81ӣ��{�V�[&%�$�ElM\��y�!� �i���_��ZrWϣ�f���d�;�~���&���c����&�re@2���C�3"�2�,��h�@W#pbe4��#�N�@��~���"��":`�����|�\���ȏR
>0��d���!�9�84ڸ�r)MR�	� �.5y$��Q��+e]#�5"<��������J�K0�:=�P��ba`��y�a	n*���}��׾�J����$v[z~�ϳ��dgT�T���C�8^�V�*��D��ClP�U���b��a������$[RMic�4G����^�2��-����U_曡#$�����=��dЮF�Ys�x%.E($9f��B�$@���! ����tm^j�ԣU	mb�AD4L_�F6��"eE������(P�����#��B�dB�CL�RJ��,�i��4��S�W=�v1�'��.}�!C�AmA/����B�|^ڼ�䂴�!j�\$B�slZr�dX���%��P��K�Kލְ���p~�^�>�
ʔ���?nD��KF�]�����Eh��m]$�I�V�-*�H*٣9�0ho��٬H�@B�h�R��ԉK�	q��/o�$<�&��܆��>�;��	�,r?�_K���.���DC)�H����@H�&� ^EN��١�~!��1x@È� z��̓���O%_����ɰ�����4�$
������	�U	�+�? ]��~����Vj��V���]��|����N�kg�6i(�Np�3�m�;?	�O�dW��z�2G`�G�fϳ�.���w���X$�~��3�}�!��W�00B��d�q����'*�:���h�����͸i���Ҁ��%�P��(�J
ĕebj(�%V�JkM�c+2u���*aX�>Ls��u{�0���P?��H����>�����="F̏��
){�� ��3m[gY�"(�еiQ%����\c"
�p|/�4R,XR7F��4y
�&���.*9 ;�w�#�^�ƿw�^|�n �����p�L����5�PH��8�Ƞ�{G�����+d@�7���GY���\� &�J-�j�B1��d�`�ڎ@��,M
��!����Md�!�E`�G�X���w H����+W�߾@�����| h����^�JƵ�EV5�
X�7�-GI���Ĵ4R�����=%*6nRd��!�z2�v�p8�UNV7BILpE�Z=fK	Q�a�h2��K	"X4�x"�;��0 �)z��U(�5�N7x	֓Ȱe���<Ȏo���b����4��'+瞐I?XOG�W�{r ��H������R�v� ��K������VS�'�M�0�ן���'�F���y+�_��y^H41��@���������>���]�=i(���M����w��,�� XX�i�Ql�F�".*��O��e���p�}�� YU�#O�����pzB�~H
�ސ#?��=h��([��%"'�3��,��>%Pڮr)J��ꅦ]����*� ��i���#HB1�O�O�[�{�X��-N�����D����?�J'�G��H��3���螱����q�a(��`�#�[�E�K�����l��k\8�+Q`ZIУ\A�ڷl��h9���Cx�)���/�r�<_��q���q�k{'�M��O��^�=3�Q�O�>��/��$M���|�����]|��¼���W�>SJ'��r���Ǫ�#=^/<F#��SA�� H�)�#6�;R�a&"�[2%;ؕ��k�_��Ҋ�AH��bg�G�8�49���+�^p&����M����T>�B���"�}XV� �4�o�؁������e��B#��W��<�?�#��Z>ޕG�4;�x�_�B�Ax�����K�?�V������'�F����f;�P��fE��,�ַ-À�]@1�gT^	I�>���k��]�G%疐��1ő�0�,���*Xǲ�u�
��ر�L�" E)}+�L��a��N}J�	 o���][���A ��zx����?Oѷ�.����'>��'�7MC�|���L}�~�b>|�\H��D���I���Y��{^ְ�6iR��8:�&%�l�A23���@��@�X�!7hT����q�BE�j�bّ0֮�$"��(փ"X�F�7�� �@1��@�����x�+���D��	�*��2���#�� ^��#Շ� �btB��F~??��	�|�=-����|��=�H&���>4�:�z��#���I��$� &�$�L���0�n,(����Q������h��H'����^������B���?4h�f�a͗���Dr#����~c�>I�����=O�1�~��V��$��F�K6d\�X���R)i>�	>����:N�?s��N| ~?��|?~�3� �G��W��Z4�?��i��6Y�p��'P�ʚ6�)k5N.-}Z�%p����^����r�s X�kd�	2EŌ�3�1�K'B�v5E�7}���p�\
WRA[&�x$�=᱖%��+�h�3ʓ��f*K �h8DL�Hc�3 �A,��q� �D���!��Ä�� �x�J�P\�.���$i����2�v,$@$A%� ҂�D\ٛ�X�kBIc� BK28��ڠB-�^!H�<�уK�$��J"�G��ѿC�|	>w��ւA,&TŢ�E�Ђ��Ř"�@��[A���W�j��� �D��M.y�'�c� �_px~a�|�>p߫_�y����8��g��<7X(�!����#�ߎ3e���������mI-j��lf�fe'%��v�P2D����8`�����ԣiO��Q,�C��Y� �|$�	0.��?k��X/�����{�	'�8!s���E6��jR�j]��A#JC)ՇD�X�F)�mA������KKkY��j�Vk!r���I�A�_�{���Y>e���n���j�<*bX�Q��e�O �b8RK)��!;�*�V<�o�bHD��a$��`f<O���B �i݁$|�C~��	�Kd"N������,e��ۂ�,cdŝ�*�hiPH�0�Y�@��
h�c��b�ΐG!�$��B�����#�{�d`���5XHt/)X���,vh���42X�p�o�BM���96�(zT��B,�TH �`�"�Dӊg&
�&��Qw�.#&Ǡ$�
6O�d�2�C�n\A-��C��o��W��D�g|��c�
	'+Na�R�-H��,,|��9���zNL�|�� ��I�Y���A3���/<����J��PH,�$L�"���
\�7Dc�$0$@U@����"�%����`��i�r`��N���J�S	��VL0Ϭdd�)$���i�٠ ��B��I�$�~lV����?��� ��?�����4e������GI�oK�Z���3@��Mn�R��n�xdI$Jm�%5(�H�M�:Y�RCW.2]��\dd?[�%w��f{�S����>jC��u���|j�t��#!��I�9��F|'2�0%��aBф�����?�� �$v	$}��?c�`"��B �.B0_�����3��=\@�.�3'�|���@7�����G���cA>0�B(xOy	�NqI4�P�j�����%����("�b���&�K(t Q���"��� &I�Aq(o�� �Pe*I�a�&ԋ�T|A%����$��K(l�فd`��q!�	�n1��@A%��M��K}w�pA?G�����{(�!띛�͉3(0�!܁i��2^a1��ϻ�H�l���x� ��@ZI���($CN�3�g��h�Œ��nn���bte���Ȅ'٩���Y��~BȀO�9���jBa�"&P��k����: �bX(H8�N"��@�(�)������6�0~%�� @��O�I!b	�	I$Gҟ�|�����h0?���8A� ���K��~�x�1ACP�Fg�.'��ϑ���/�L��'����%b��%�,����C�)M������MŨ��&�Ay�b�A�,��D�~� I�����~�A�IA'�O�ϕ#-:E�> �� ��>�#�N �D���W(�?
4	)"
#���Gٲ(#�`딁?�s�r|���L�_S�V�_ʕ���*���(S%�-	���U���H!�W�E�}��/�6{>�?|��U	
O���������6n/�,���'�x5Y�>������B}�� ��+������ϙJ_�~{L�r�"C�h( �D��4_K��Ա3�����H�?���e�G�u��a9*��./���,��`��)�Y�$�"�X AX1DF
�X�P�B�Df�/�ꑗ;�$�·u�ƒ�w(��ռն���{�R������	JB"k$�3��������������
f�Y ��b�"$E", $ "'P����@�
�_�~��0BE�0�14�8�tf-y���s�*�V�(!ς�v�/z��I
M�#�w�u�ʛҦ���⡰�<��,ЀPb��侙
�@h��"Kݼ�~%.Z`�T��������~_OĜ�3@M�f�@3��d��*D�����z>3���?kǹ�&h4
(P�1 �*A*EX�RA@�{�iDcs��'9��߇���J&P�L}��Z ��Z5�i���#���ݙA@9�% �H@#`��79Ͻ����A�ː�HX��I���vu��jE&��3�y���&��6�2IL"h�0Ebi��BuOmj��g�Wm�#	����'!^�[���̠e�("�B�" @P�CukY�Z�hh�WU��'s���Po�#J .J��''m��;o�E�ȱRAY]Ã�W3�8�]T��# �t��^�'Y����@1D9X��E��g��8ng��R����O���$�I �B"�)jk�_U�S�LJlq��9�~��=1�8�����ixo��b���xN���0���:g�X!=����7"�����OD~4K�hr�	�\�����4ij!��>mo.���Y�w�[����t\�ɇ�������]�
cb ���:���Irg��?�~~���{|+�>`������w�C��=}��X�rg�(���O�r�8 9��"� r�k8n���m��ȆC�}S�2ÿ��z�)��>`��>�9W��yR��Ec�i(�Q�IV��lX�Y�F�Q��_�~G�_�U_51��MUP ~>\��>��]���d��)�/��gt��a���l�*���O�z)�C���>_|F���.�����R��U�EABEQaى��0$dbO�WR��DcY��T��&��k���� ��9ĝwM9]&s��n���h4FM�6
�[j"M F��Q"(�,#m���:���ǒ�	7YV$�j���͉�$IT���I/�ɒfd��>��b�U
���@�o`OX�JB�L>�s�l�Tb��@z��V� 	�WGd꒝'ѓ2I�&N��rH���y���n����x����J�t�7��y.��w�y[{���V�ɾ:���X�Ţ���h�J�
��R���ct�EP�����v-�lt1�� i�������W��.k��S���Lmk�ί:��Nr���ѓ9�]���w:�)�]wQnÔ1�wqI�6D�\���ZI*X��;�J��_+������������{����gkS���#l���m�6[�D���v�Ͷ�W:�6����+G!)X*dqp�0�x�HX�8�1 ����-T�m
�Q$J3SB�:�6���
�iZb(�C�P�TALu0����
�	UR���U*Х"l������nK'x �b�B �P !�	L�ԑ��U�9.�r���3�298�}ݒ|�8��ڒ�Q����f�@�|��HE���"�L��3�|s"�$����V4�P9�<�L�Aˑ4�C��ԀNj��]d�-�LUd�����{>����XG��t�ɂh����;��t4E���i�H���l��lU�{33 G� K�,��P�PVX�M���b�W ���������(:ȶ3.-!�!H^\8���/�bO��^$�!,�0Vj%
�K�!X輁t�c-��Ŭ�2��v�d���-y���e�K#��#>f
���ǌ�`HXI�e���&�˘�<������d�!�7g��rRG���#<cO���=}����ђ�y������^QA3�.
\�ͲTd1����gfR��L�-@.�f;!�.ax�^!��}&d���zo��gdd��n9��HşSg��$0�"��4��mX@X�&ϣ͌$��I��]aD>�!c$IE��c�[B]��R�,�܍�U�K &�5ɛ\���L�(�L�RPY�b�B2�$��(����h@�s�t��
L�Qt$$*J4QA�qau\�J �R�K-�����X������ə�}"zw���'Ca5�����	�ܲ_��\�Lo�{��$��
��"	 ��Ż. -���Ѿ嶌�0�͉�(�(��X��5�R�ɤ&����\$��	�T��Ă�`��/TAI������&�t�HB}3�>�)���"�Yd\Z!�U@�ŭ��>
����� q�
��Ptj�ۦ��������$� >�n���?c�������|�P��$@#>�mkM���_��}��t$ �H�*(��H
�v�y��UJ���5iKl�ET"�;���c��R�����N|�Ƙ�FC3�S�ބ/�_A$DaI=��?7=�1):U�Cy��Oۗ�l�S�?���I�bJ(�D�c,�E��>������A��8|���#�`��̠c,�bHcA�!��0���]�V�"�@�$.H��V}��	�-�K�8OV�UDȏ��'1,h�w�K�3�4���p���ߌ�}��4���܂∄�� "?��u�-xz$����S;�{��||x?opV��?IX���A�?)��o��\������i�I-׾�����bmI�b���qc6��Z�tǰ����:��k%Ү��[��r�j�:J!�c
ŊG2�Xhђd�vl��{УN?l����>�7��>��2R$�d��A�\��?��ӽ�|��bq-�����d�|���*�o�&4���;��@����Vas�/��7-��g�>,RRB�xNDB\���ơw�a�HD��]�)?�!�=�v|9�d�!��~� ���J>/���>��Q��M~&<9���??�}��2hG&Ȅ�=)��~K�2E��R|��̊(�ā��P.@x�
��t)N���>#�f���B�|��O����	�xی@�j1 $$	@�|�Ct"�	�/~�e��Wz�g,Vb�M#��}���(q'	��N��c8b��'��X5cHB��Y͏e�P( �*���b�C�B��=#��u��ܘ��POpC���ؑ��(~��>`�^?s�p�xf �����ƛ ��ݠ�}ȸ3�$���(� ��*��^w���y�T)p ��T�-�� (w�֜'2���P�:���7�;J�_�(���
� y��"�A��pP8�	w���]����|�L;��{�ཤנ
i+��6�~"�⡄
F�S��f����V�Z�+j-T_��m���&4H�6�{+'G���������a���3��;w��A�?�;?;J%�D� ��)�y_5x]�|3dz���>� ��m�i�龑H�tEP���>��0�D�?o��7 �F��D~a[}�f�ˮ���m�mM$�D�j��ekeZ�)��L`T.�bS��*q��';�/:��v�{[ikW�I0D ���XZ&b�@����	J�n���J(�K��( @@���] ��b� r�(�`�����1���"V�7�|j���Wƥ�ר� ���� Y# �
,�)����iV^��m\K�/!�Kk]�������
A\S��LUUu�CT(�������EH�L��u�!.$R�q١##TYQM��!����Z��DD�$YQ��'=Y����j,X�U�{3M�v$LB.�y0Q�N\ِA~�î4�C��:�J%�c�� ��GC51��5�h�p�q2��^� d��flJW&$�<ꢠ��˨��J;3�ߴL����J4��\����4�>�7�݌�R�D�BI ~�q:��@�l`���\�"�bE\j.j���6#	��~�!d��&k�B����-Ujߝ����w�����`8��)��w܎���M��0x�\��M�
4AGl8�G!j� �D�BJ�>USPl#�(ƨ�B"�^ �!;�e��9�A�7�� �A1 ��GP	�����/.)L{oݣ�|���I�5Bo)�LP(��5)�

��+���%��	�C@�� 4PUD�?f�� 4r��DB����u�3xts�*`9D�3 &1����� &Q#Y��3 `�u��@l�`n[��ڭMje��Z�F����d@87��l���(�f�⦐�t2x4��� l�	���L��f( �0sDŀ�mGby�Q8�s�ٱ�E�w��w؍�"c�'Ż���kE�BH����v�q�����v�UHUUJ�7%�t"2 �xb�٭�J"�� ���L�eě��xx�>�dEdɌډ�ė&�<��F��Uۄa��H,� ��]��;��ڹ�
�I�].;��PV60Wr���7k(I!�$���q g%f�k�v9�MD�:�za���!L� b��P(кN|�K�a	BI5��L ���I"�7Ŕ��F��M@ ͚���ij���F�C*%�x�1���(��'�A�K�!���A�;}�f�`�� ��vFq�����i��6AYXb3���<Nq�K�At��v#d��<�Lq8�r�ub�!�QP�Wl�qvp� ��ɻ2�PnCI;jf�b �� ��E1�7^މI�l*э��)���d1����5PʑN(�������(�S5B��!���B����ʆ�H�Cfk��,8���u�C�*�C����s%9�UX�Hڙ-0LW!z�y�4�(T���(C.D0�)"�(XX�P��*�Y��QPM(���h ��p�(��+` ���H2�e��"`�Q� ��Ǝ�ӹU���C���\d�P�8	��*13 �@t@ӽ��PC���p���(0s�\9� b@�x� �%�y�Jq�&�C���&\�xGUU1�^|������ �>����e��`��01U[V�[��߈��jlTEMEP/ 5�p��އ$-�.
pAy�)�n0G7�:�{M�h�2���f۞��׍F(�&ϔ��~/T��w�M|Ca4��T7;�Q1 ��Q1!���q��@ 2C^` `�n�D D
".��� �Р�cr�d�RL��㵾K��9��/�bG��r_��B5� pn=AV�M0X  �`T"�:�5`ʭʩ 0L�g��.A�9���4���dr��Sr[4`'� �D�ʒ�c���aSn�!*���0�au��� i�P !ď��dzQ�v�<�����%@44���r!�����u�� ���ِ�!`L�1��(�78r����rD��P3�AU ��6H�ZS��b,4�dϠ��(�d@�t#@�9��頇 �= � 1|v��H )��*����]��~��tLC�;��)�;�C�@���bpE���!a� j�m�p.�9�&�fđ�e\�7Ⱥ#�r�j& Q��32rϵ}�`7�}�f���$@a�p���ዴr[��d#}� �kD�Q,�����^+$�� �\МME�E� ��lh]���Β>��z3;�hR'�������^EA@�Y�׊���{zЇh8ԥN��9|�8������Gw�,hw ��1P.}��~K������ʀ�X2(������ݵ�HB/~ }����u��B7A $$DFC������x~��k�0�<%�-�^������"�^	�dD	Ӵ+����N����4�3��`	����� %�;��
H���BvX�?�Ki�o+��9e�yC�I�ò��x��}/��~����O�2f����9��?.��3������󶷝�����ry�s�G�w
Uq]�p�
G��r����'5y]�}�H�Z �+'�N�ӏ~R�_Җ��dKw�������	 ��JC��]wm߂Ie9�ʐX��ZȪ�"c��h}�Q �;^�K� D���?�Б�K��*� �϶��XG��==j����J�tq�����M8^#Bڹ�S��nC�yN���o2�G�{����y��c_�_�שn9/ݵ?gǿ�����������a�o��B���>�4�����Ч�ԏ��,� C�/�i�� ��y�e����B�?\>�pl�AGa�w����M����b�_��yn���������w�Y�����c�����������O���K��~�D�O�����R���A{�Q�:��A���I��G�؆����;���O����Ȉ���]��s���]x��ٓ<i�x�'�/���h~MG�S��)��'��Tg�S��~��~��Ǡ��?�K�x���_?��o��L�gY��j�'�ڗߏ�C���}��_�jI}���������g�/��ꋸ��@|���+ٓF}����?_�=�����M5� �������wk���}o��|�w-�w�=w1o��8��������]v�Y>W���l���wNc�����������ݟ���/���{~S������+m��߁���������Ձs�d{`4�$��t������B�#���]:�������r��O������;���~���cڷ�X��⻖���u\gz�sH(~(�H�줛b��:�'���
�@8����G۷/��N�������u����m�f�g��ϝ���n���]�e��;���ߏ�o����������bͤ�QS����?9������������?3�)��_�-����_��!�W�������\c�F� �v�/�����������=�����~)=�>�I	��������'�.�I��`���;���������y'���=G������%?��Id��^���|I����?����������������>��_�־G��}g��_���W���D}_�+�e������l����{�#�~2�������ϭ�)#i~o��>�w������������hW�1�>����4��Ȭ?���ׇ�����1|o�����Z@�ޝ�c_~���$�����e7��O��g>g?_���ߟ.#�Ӎ|��{�Q�	�����}�ū쾻�����+��/��_�=������#�?-�M����?�_����*�y��~��/�$?c>��l����?��_���Y���f}��}_�}/���������}?��������i�_���}����V狼�<�w��6�N��^[�����f�@K����z�'�N�����4�	#��R��*��%D=G��,����=��(������Ȱ�	�b�?�TR�Te�
~���Lb���bi3 2ְ��IbB��!Y���X�t����='����\��Q�PY�=W������$ �����\��{.}y����� ��� dTC=���'+�}RBݟݠ0����E��������?��ϙ�s����o��9������<��3��:;^�����m�]��T7P�\f~��:����9�r���~Z�<������[y���n?���y��PP���xo���99o7��'�&i�^b�HY��{�V�X�A�UId �Hx��蟟�K�/�;���,-�AN�����zR�e�"?�?f�����&	�`���H�>�Y}��Z��\(; �EEd G��~�k��������x3��y'�HK���՗��OM�߃/��𻏵�os�u�/�=�����닼~?�zO��5�[G/�zUWOF��������"?�e���	%�#��d�@P#�$p������Kվ�W�zz���u�1���_��|A�"v(;��E�ˏH�_�r��?�a��/}mB�?�{��9�?�zm���5/�c�z;b÷�d��Y�x)W�� ��D�+=�L�"サD��EϦ��	ƃY �����:��j���*��!�b���~(5]@�K��+�r}	J���hCq��6l���,A��Y�#�Ϝ��l:/���K��� �"e:���$�u�~a(B�w�
��7?G���7���Ъ8� <g��>���/59H`�C�yɜk�I!RQ%|P�&B����_���ǡ�0�2Qx8EBAUx��È�0�a�P�`<���M�+o�9�C�������u�{t.|����(�dO��-�����}mEl[TV����$(����H�Y ��HB���-�ġ<O�%}o��a$�X;�BP"��"y�����au�ϲ}Ą$��PK����#�������`����A��~�������C�ǚb�I����a"s&�F��`�����D��r����]�$(�FA�PXA y��ˋ� 	`��������)�H�V�[���O�8��!�7�ǯ;RlC�\X�>} ͷ�O���!��e_�}���	�������1R(�F ��*�,� �=Mu�r#DU���\�Q��EU����YDmB�
-#cM
A(��JT���Q�A�$D���������H�t�@J�)B�
@*'d�(�� ,�>��$da�����AC���o-���R�-Sj���mDD"�U���1P���@dZA,)R�A���V��>Ӯ�u�u;����wI�nj�uѝo�g�|���X�:�W:H22���ԪrݖՅ5oK�}�z�wFSH��w�弾���}ow��ș�]���ǟx�h u�)�I��κbW�Օ�S�B����UaĈ/T*�D$EF�����F�����-<���j�`��a_*���j7Hε04��N	ʼ�x%�C��f2rbGq�t�V���$�֠0H�s\�;"�[ɮQU]u9���P��L�@ȉic�dElŁ�A6t驊�=���ɘ�ʬS�d�&w��ٸEH�D,�u�Z�Tښ��[ei�KR�5R�5ek+JҼ< y�����ď���w/����:w�/�n_���m7��,��9Ic<^�KId�m]+ږ��7�]�,�}���B��ԫ���W�5��˃_U���j���(|���"$O��}Z�nd6	=�K�?_$�uTO��~�{?g���X���;ߐ~���_h1���=�u���_W�~硗�R~�u.��w�")��s���k��є�\Z2�n%iN4!mw���饩��J��5yq�ύI��(U�3�2!"�`C�+�1M5t�c�~h�z�6�$���
�Rb�m`���Vْ�o!�U���vI�Z\�L�zN![#;�+IN5��s3G�.t�,q�Rѐ�%5�^�\�<��'%Q{��r��\L��啒�^�A��Q�Z�uk��!8?3�������pl^���*�IJ-�Wષ�w�yb�����nQWI��f|p��Y���eS(�e$��qz��2�2�5����ۚ�r�F%#d|�k�i`�,1��m*l�� ����,�a�V�a\W'ր�r���A�*a:+�\)B� 2l�� ���$�$�HH"�Y�O����1ߩ1[5�]"�X��qze����3�Z�}��2�/���2�t�~�3v�ع��0��H�_:ʶ�����K���mvhjչ@7{����F�`�Z�c<������\�8筶�_Z�Io�1}p����:oʙ�7�Q%lsʷ��x51m%�2�?:�lr'`��xڶ�M"�t���?f�5��#Km*�����J�,v�E9?]��:J��ع��+I�;Ga�6���vH���"+�[��o���z絞��Q�W\"����W��%�a�5�N�Y��yK{>��5�"�I�TK6�<tW.�?y�|��m���)���3�]��[g����iJ;h]����_�T��g�D!#$!B�@AR@�0"�[[Wq�����q��߄6'�]�� ������GK�}7��'�o�{p䷛�lW�z&s���p�0X�\���-�xeL:�P��4�myu�pˏ;�9+F6�$u}��^Q�8�Ә~�nV.�b8��[e��b�b��oλ�vɲ��Q�,-}ߴ��C�A�[�F���zo�n�JӌyW��U�P�F��x��xC�������;g����~H��wۚ"��+��x��L�[�٭�:VQm�'��;g,��|u� %�<�W�s��6�����G^��Sۜ�����~ϕvкvq�H����q�-<�~�t��,�2ˍp�c���?=�[xo�'\٧|3��LkkSka|W>mNX��NBӧ&��>�-3�����VӔ[Gq�#{O�52l"�3<���X�:@]��,růx~��8;���oʹ�U�����**H X� �|T�F:r�Q���ƙb0���60Y$̴EHX���`�A��5W��U-�[*�jj�jVʩ�(� #b ii��s�+���MM�V�v��]?����ih๽ݗ�׎��7q���5��m7ZQ�Q�:�1�#5��}j�pˇ�
`�s0�7�:�m~W��ᳫ��!���:Q��ˡ�ںþ��
$yR6���F�ݫ�=a�)Tz�me��q��`�'���4�}�0�>R����}��ќ��Z��;���WZ��o���^�B}�U�v�<�$�F�)��'t�n�ʻ��nsƖ�k��˯�5��&�W��}�kx޶�3�y��p�WJ>�7;Z]m�rҗ�b:B������vl{G���μ��<6�}uL��m�\ڒoXCs�ZCN��چ��	�(��?)H_3�^{���.���J�t������8t����Xi�[�qǻ[ۊ�}���e8��~��h�Xpz�m}/ǥ��9�ݻ�dv���4z�t���|\���+;���~�>}K�']����r[s�e�|{�S��]3�]�|�[�;S��u�P�u�t�� k�n��9�Q1�����_l캚��*�e��������QB��db%A��_t����l5~�&���3]���B饾��]��ڔ��Q��9Z���x����k��[����S]�t��O�}'�t��̝�i�n��~6u��N���Ǭҫ�<���^n��ɯHg���))�^���!�zE�PL�En���o<+q����|�q�����w|J���;zE��m�>�����z���RÝOG��}+:���t��6�k����]���O-�?]��>��}=a��?^��3��{���ƱǗ>}W�NY�-_OMF����?9禎�}2�Ιr��׌i.yέ~r��8�K[��u�GyǴ��k-���hz��q]_篟8R�l;ْ�M��b�:R�P�ij��� �^���@g�ϛ�jï1����_�;<�t������]1��״:�:jg�7���8ǟOE�>��ꝫoKx��������-ӷ�^�\�w�$#���w˽;Tp��˛x.Zs�<�NVDoq�H��Y���+Ӄ;����H��q�%�������x�/_7�iY�yӽ<3^���{��w6��}6��<:��;=��]c��w���L��|�x��=�쭋��5�x����+�ط���a�N�5�_^��9�.}_Ɨy�l7���tӈ�ҋF�~��0c�1�e=U�`� 0Q� �iɡ���4��{��m1n���;���[�;�N\9�8��E��1�xM����o9N�>޺;���Y�m���|�V��*���� ����}<{D��m�4O=J���Ȣ�c�z���DN����<% ��?_9k�}*�;����N;�>ޚ��V�պQ����g�b��K�qĴRl�3��S��$�E1�� �9"���	P�<[#=�$���1*b�;�.��B\�J�g3�	S�!�N7C5��5��u����$Va�a9��y	g5r�ed�XV	)&W%8^1��NX[� �ʉ��iu�U��j�I��ľ<�_�|y|�X;ol=����뭳_:'�"]��n���W߿�F�wN�ӛ獛l(Y�u�s�zD�Y��4d��e�2�MtTh
��c#����s�<#��/��\%�\O�zv��_���{�����S��==9OOxy��w��\:r��t����폶{M7뢅\t�i"8`z����z�I?�
d=d8���_�\-5�1��\U3�>��{�6���v���f�]�^=�g�=��ѱ�=~>;i���Hq��,����K�K��A��M�5�R��nǭW-��Zx�~�=���|1	mg��lvww����m��|?����0��͏ŝ��
zG�;����xU���k_��L����ͭ=��73g��g�\h��uP�n��n\�c�v�q�����p��E��VZEF(
V�С�FD�Q�m�(��O��{���{c��z�-�����1p���\=~����h�O�8D�Ҩ��Q�2�[���_�*i���L#J5�k�ې�Ǥ�7���<���i~����[�F��������#�6cHML�2�J�E#+� �h
%�:ˬQL� �Gl��i� %J��	�Ȟ�r�3�a�� W���ea����:l�<`r��m�FW����"��LqE9VP���h�T��%�b�T��M��i��Q�	} �!g2t�*\�a:��H��@Q��'$B�+m���X�	mٟB�)\œc'qX�mTT:��V��'�H���k�t��1+%..�\�ۏ7��:�?Y}�;p�أ��V�[\�߉�Ҿ��g�}�̙y7'gG��H5�����xy����6��:`����=
Y��)�e�x�(�5Yf�Ĩ�1o8{��=�s���-ۼ����x��{��8C����w�K��aW��W��B2lhS��A�zL��ϤK�/S��TB�.�M$�渍C�C�Jf�hI��2Т�&C��k
;V�e�������z�F���*;�F�T�놺|�d�xj�2�)�� �m�+�)C�Y2�"�Qc0��d��$VkƑ$} ��)�jPZ�vI��}9�-`<느@E�c�F�I
���XWb�k���؎lԀ� ��@#���ϒQB�^����z���7�aۯ�0�Wս��b1���y�O�^xf�˵]P5AH����()���Mi��R�j�T��H��E"""�fn��
�hzA[vQ�!q�	  `ĥ$#a_�[XcUdH�V�ꔅ_{�G��~�:wㄯ��o����1��N��O��V��Q�a�4�B
�� ��da��f�)$\	�p�=k���0h@rd�X4����H�RHZ�^_	y١9�!���ӎæV��B���JĞ:8�7�� �B����d�ZAt� �5x��͠��P�*6s'D���鳫��*��H�$�;5�4�r�I�@ĠU�m&@�e1Yr�c�;.�a��"�d$RD�hP��Rb^V�YƯ�5�\C���Z�C�LF �֜��	�0��ʕr'={_^�$q�e�*�{�=eF	B�"{�[¹�]�.4q�Mb%7� a�7C:���Omև�x���b�!)�`��2,$�l]b�M��(�iXD��H�g<'dT"� bM�B�AUu�y�^�Ё��r ������}�}>��8�]��pz��&��%dot�^��;�xg+\���'!��Hp5Ņ��Ya����c�u�L8TaA30��4�A7dq�`�B�II1m�t���C��߂���`���n���Z<�����9��o��/�����<�v	%�	Q�j`WȥU�8�~��"�B�!e���%W@��Jo�~��魻e�^����a�L��'5��n��ˡhx�I:��v���䍂TF�u;Xu�ݼ�ᐒ)��aș�0�P��:}RZ��T��I�����0�AL�abL}�H�2��$���[�j�k��X��E��Y���O��SX4l��@��=p�%T0� ���7L��!$(��ڊ��p���SYD��`wH�\x�^[�aV4i2^p*��.� 2dƾ�L�s�O���?��㵼�O�����^�ǰ� ` ��c� `c��1���c�����:7�oE��=rD3�D����0VL��k��鿶Q�}4e��E�%Ǻs	�4('�{T���QBm�$���PD�dQ_A�.���u5��
"�[�(a=�IE�k�g�h���wѕ�v\$J6��甩�c����ϰڢ��w �ae�ZT�e�,��!�dU�7 NO�)�-��1�#H��E�dlRF<��f[%[*M)�9�%�$��h�g���`�-�Į����]�))Ap���L1SA-*��"tB�k^.)(���h8`P��XLQJ�Q���@� ���$y����b�H�O�Jv�ݣBy+t�@{� g��cRT�V,�S�8kI�q�g��eB�״KX���!v���	��0+4�1����1r�l��"D�ȋ�$�O�i�CԭqΦ�\��*D8�L:g�VCW�P0�
�A鮱a�δcT8��P�j�5~�o7Z�Gڜv�͐���)|�p�'��:�"V�`7�R�`'6��ةuH�4��q�\�ȴz�H6�	��LO�h���.=Ha���I�I`�Z�� �c��޾�9 �s����Z����|�gӍ�ze_�:m�'(�&�`���~I��nfD�Jxn�
�:���A�cP0i��'.b,�=���$O�+ъ�(vTG\������6Z=�M�l�M����ml�2m6���� ��"c%ey�����R�]g�M�SŶ�7�9�B@	2贠:qk�|'�㣩"$��OLQ�爉�D����E�|��qY��m�{��8�����ڋ�D�Β�FNs�,��ea�^v�'��� s�u�\<7�VC��Qx��c)����>U���*]���1W��U�B�83�AQle�5(��@�uy�	.�[ɒ�o�����Ai
���Kg3�� �Jj��jh5����W�A'`�d�����߉�:��T]�P��p���jn@Q2)H6x
�	4v�]v��U��(!����$��Ek���<��9�uk�&P����6���]Fa�e�/���:^��j2$�-�B��Q�bm*���Ҝd�)�1��Z"�v�;�z�y	�M�$#�A��7�d�WQ�ILا���j��G�}��eK�d-X�1�FYm�E
\/2�4\�%N�kEZ�GӵS�:�Qz�b��1�� �K*f��B�;���I�hh��{ӵ�$��`*f��yA�͢Bv�(^��Zf2��׃�0�LQ�-� (������U�<5+�D�����R�lP�2 �P�3RC�묲-BԱS�?B�6���O�%�ӈ��J&�&�"�̛x��pA.@�"y��m�1"���6[�^>�<�@a�2L"�`�NYt��NS3�d�
�nefU*�b�3�d��o{�_YX�v6/MmUT�)�B#7#lT񆥅��p0���
˷J�"�R�`j	�5ˮ�2u�k�9 �8�ݜE�4�Z�i4B^��(���3w���J:��F���D��ɶ �K=��q��)#��H4qWA|t�>Bn��1��H|��7%&|̲a�j�
r�c��$s�	Q2@`��'NR��"�E8\սR�M0íd�[J.�����a%]Eg<��2�N6��Ӎ��f>�U�LONL�S^����,Qo������>�E4j�R�K��옯(o�Ņ*���Z	��
ɉ� ��Z�	��T���F�A���z�l:Z�!|V�k"ﱻ�-���L �]����M��`[��Z`z%��бjؐw�2浸`��C,�L:e%-6�k4� ��Z"��ƕ������㶇�to�\�N��?�(��C���f���e�	�0y˲�u�M������y�t�*����;�\�����hg���#�4r-�@5Q*c��]�a@`�>�`�Pp�
�vBԪ%�Bcu�#D�����Y+L�Oh�դh��3�3`�e %Z�h6zþ!�C���5�d�{�o��7�M޻s��ux��~���o�S���w�-���.����5��������^��l�*۹�j�?f���/�?1滷j���ܷ+��R�")iVJ�!@QH�J����^^"�Sm��K`*	��,I &Ys8mZ�V�m[p�Q���˧v�F��Z�^KE��UͶ�-x���y���r+-R	)F�JaD�k���6�,�#�#��� &@��)�ƬlZ*6f�51[6�(׍ʍ�EQ�э�h��Ʒ4U���j*-�A"��hDHA��e�>o}��~_�}�E�>�������_�����d������������c����W�O��~�����������
��������Ș���lR�W�_g���~O����y���_��V�W�~ÿ����{��~��T����ȂeO�`_��Y���]`�z�Y���r_s��r��O��<ߗz	Nx�$�	$$����lEcPP�L��&��F�Ƴ[kF�h6���Z��[V�B��iZ������Y$�E��l[3!F�&�T��"(H* �� ��j���Q��ț��j(�("@���H�m��kE�ƵѵEkF������mX�jѫF�V��Ub�Em�V�km�jڃUX�Z*-�����[m�j�j���ڱU��mU�kh�ƫb�ت�-��[X����Ʊb0X�|Qap���k�n5T[��/"����׭��?����������?�Ke�~�����~/�y�\������?������{>�z���}�>C/z������=����/��p96�~o���~������|?{��������[������ӿ�򿉷���������?���������o���G������{n��p�G�p>3�n3��c�����}��7/�����z�;�|�f������x/M����E�~��}����e����AX�|���U(|�-{|����H)�D��L�l�3i�2�H���L���1��C#BYF`���`LQ�,j$iIi�!(�(��B�i��� �L��)4̈�&S%D�$�1��CDR! Rc	�	��a��3B� �0L�!%0���If#4(�DЂ4��H�4�L�d!���(С�
Jؔ�#"34&H�$�0��2�i,2�Ta�H�1�d4l%$������6&�4�Ld
jjH$)D	�JՖ�(���������#������}���z?��|N3�=�����?���^q�>�{�������.���/��~��=����G��)x�ؖ�D��������jux��u���=_��?s��~G���=�{�;����[�|ׇ��#���#����wO��6���u�����y�쿿���s�vyس��AEO��7�;�{弧��Z�k���oM7]_��\�o\��=^���~BvZZz�ٗ�Y���-L�B��u���P�?�Z�i��q1�K�����[����-?��X���jg޹�d����.T*g���	0��q��/�"i���LO?���1JC�eY+һ�wz`�ĴVR�,xF§�}o����=���&N��F�������ӑM��3<=IÒ&r�Z��+�
э��p)#b��=C�>5R��:J�R�
����K7�!�V,^���y8�iX����5h��](��-�q�G+(�kt�`f
�a�,��٦%�>\�z7i��0Q��(#�G��аG�O�z��{�ҾP�GI�0�z�e�	x�)a�-���pFkq�����T>�NL�eXe7���: �O�G*�Ѵ�ON2���gG�]�l�ZY����r��)�i���`��jh����S	�G�a��&N���2IU6xԳ�7j�[� ���K:Z��r��B�u�OG{��P#x˼�(���s�<�N�D��[,ڎ�Ȏm�����A|X!RE�f�I�k�A�=L-	wW�E��\.���c��]Դ�4:h�3�q��F`n}x7�;��j�qk��(X��~�n�ҁ%7��������O&�J����Q)9�9�J�U���	����;zI�2k�<�8�����F�y��hpu~�.-]Á�� K:�}�,nPӄ*���i�F}^H�A��$�9�(c_Ye��U����$�G��C�_πa�m�P?A�(GfT�Fh��I�L�P�� /'�N3V��%�l����N��X'�*�MEG�![3"uMsObΝ���J��������C1���y���j'ܢ��]l־yL~�\����0B�6Xv'���HĜ��ѕ)mg�]9�aod)Q8Q��-y:�)]
����3֦ZxV5���#�XU�zcm*3f��3�VG�B-`6��ҧ�l<�~�p~��d'�}%W��G�8m�U3k�渢W̖�z�c��%�^E&�8K�{bR-�Cj�9���/(8�"�N|Y�=������W�0��\$\t�?��7 �N�U�ð��3R2��+���?�E$�p��=�k���]�K�T���g�`M�X�Q.D�İ |��G dO�<<����y��j+�>.(E
��G��0�w�[@n��\�	/�����f�<�|9���������2��a|��0�D
 �|�ˀux	�]IP$�o��.X!�j]$m�	tE*)kO�d� .��a
��f!E� �<�� O�y5羠 �AX#�Ђ!�C�T�מ
D/����<�'��.�_�~xAJ���9h_�b�����8�Q2�̚|̐�)�?���2{P�AAs�'�f<���gn��@	>�`��4ֶ�ڛW��s*�i���QQ�b 2 �dQ� L"
� ��PIE�PA�T���h�� ED�E�**�Q�cUQ�V+kZ�B�2"��ltYV-�����n�PqC2_,B�l-:!P�b�)�hTD��������Lr����]-�v�g�|.�h�>b|,�$	'���D�I� ��a-�7@/�P� _D΀�*:L,�j2��%��Pb�%�BC$ �P���-��,/� ��V(�DřA�[B��t1B�/�D*,[�|2J��E8T;l<�n.�[�]������I��t�̛]f�*ԛ���e5�13�[g�����������������|����������w�������"/� 0                                �    (     �	      3��    "       ` �     @           `5 tb�������I�      �I�R$C�    q!"EUT(�
�RJ)H�!$$H���H�	IU�Q�       �(�       d ( �        +IQIg�       �R��|   w�      � P+^     mp       0R���      � +�                                                                      >n�       ` 3�       �9�� 3��77K��(�iAѠ   �                      �@�@�    v�� �  �        �            tP��P ��        � �C������B� ���: � h Q �J�UH�  �    �       3��D       ����      
T& �44�i�&�&�����@�  2  �  CG��jy�� �M@��� hi�z�M6T�"1M         �h    ��h�������6�z0&&&��&� L�10 ���	�0�0	��!���A�L��)T�G��`h  M0      �             ` J~�$@L�&��4h  �h �   @h              ��&B&&�D�!�h2`M�Cɦ��L��L�Mȍ���##�Ph�OSh���OP�ОS�i�!��M���`��f���c#� � �/���wW�,� >��C_$@�D`�� ^�^x�7��0p<J)�*� �~O�UJ@�!�����~��.����/b�� v����T�7 8�����{�y"��B���*mĵ�eTf3!�T"0G��1 "v@p�3���UFX7}o] �Z���dt��$�� s?�;)W����F
����� ����T8N�i��1T@�F JSEQt�` �BDORQ�R�������G�<� ��C�C�( jAP��{�}�<A^, �5�cH�d"A"���?S��u8�/OŞ���~{;�8��3Ox&5l\x$����X&$y"M[u�=JE�l���2>a鉫,#�j� �U�RQR�E�H`���
��^����W�~���S�_��_Q����C�	*�2
x��ʇ���v�c+/SZ���w[y����V�mKw�6O{�='��II%=>_���/�����_�����QS�y~w@1�=U���QAW`��{�߃��DW� ���t�E�G�� +����߇{o�����نI"�޸ֽ|dZ���֋`�M��,��=����VS�}Y��:��s�q�������;.o���
��@��  3��� �~Ƞ����1�T^~F�w�O�Ҩ��`��.�/g����@��(�g��O����z���w�^��qTW^�W@��|}m�uU^p�����@8x���x��۲���?�x���p@;;v4�k^�6P@;tw�  ���8��Q_0V P8�A.V
���zB���@�;:{>��y��� �UWhAW�LPxȠɔP~�8s�t���m����˲����hTWR���Uc�ŗ�n�rU�@�U�������~������<֖|F-�U�5[��Y��	8����I��䥤k|VbY.��08,`č�|�&�q!O�j �@�)EC�XJ*�oܫg��<@���|`���X�w�d��{j��?V�Y
�y�ā�3�B��y�P���t xVZ�b��d��*!'W�����(����K1ks��F���N��Ú�}hV�((ۨ}����
B*+Ֆ  �OY�[IIVRR/�ˋ����/	
ϩl� N}xH{�ޒz|�pB�QJN����'�s�WϘ	)B$p�0��2�L��G�%�gȄĸ)��3:�+̢z���v�}�%�Z��{��q"B}C�uk�խ #Bw<hs(}���Ҍ	-��ײx*�`�A_r[���쐔+��H��|�zX'�r�P���ˮ�f �H�v��7!U�)ǢC��_E�SJHA��K��Z� �k8�,�ς&���%-b�%c�{i�!c\�g�v�z/����s���HJ��x��b)͸�$!A�bՒ��6�_�}�P�C�����ѳ�N)�L�mo`��ؚkd�tSV,z�U$�:�L�݂kƗϪk�
�Q�}M���$�a�>�e"JmB+��б�{ 2�, z1J3���X�=\�>� BbY�!V��]�z_#� z�m7������78��d��|2��a9�O5�e�X�@���=���{$ %u�s{ԕ��#�,I8�����Wo-mi�Ǧ;4�����ү�c׉��qN���a�^���RIT�d����o6��곗�[��я��n�@��� �h�Ǡ���Hwm_���x�\{<�Ώ�K�m1��+S��	/]4��|1��+��@)R���0��/��k$[o��x�N,,-d��!0�9k=8@�gϚK�� G��w{u�"�̲	F���f[3HR  +ҝ�/E����>�H�@�.XO\�ʾ=�@��L5�u���qV��^�P# x�ؤ͕$ ��)�JFV`�	+	ǯ����(�Y�z��X���wn�F�y��ef��_Z�m�m�,4���W��f����c^��q=�I{�)WZ/�F��l���/Yg����<#JF�Nz�)8LQ�^{��=��)���R�}{&�n�Xz��]X����IBD!Xs6w�Oe�
�0��V>P_g���1>�L₉�o��Ֆ@!-���+�X���{�-�4�z�}ݲ�+5����Ϡ%���=	�edEEH��T�k���!H��l�liRf��)s# �'���;E�ًl�����ᬄ��QT�c���g�\Ws�a }��HH[�kN�E��K%�-�Y���_t��=v��՝�:�"�օ��wk��!I��*l��1��� �������d� C ����&bw=��0����W�-@�.��d�<k�W_[�����͜�6�8�b�$kI��p��� �4ώ���e ���px�oY(J�#�,��uˬ(u�3��|��7q�k>C�7y�[o�K�̜��빉'B@�g��=n�k��	�t%�ք}�v��wbL��.����`�bZz޺���Z0(��kU����%ib����&J��Y�0�uQ��T_�mÎ�z�8�	/%�d$ĉ�x�c"$��ڄ�,�+1fT�N���ddn�9lݽ��8�ť+�����c�{�>�Igy���Wx&�T��W�]� �cU
�����C
����"`@�Ei)6-�;8Ʃb�_R%F
����(�ǩ+�U�H�^��gs�Ab���+}�X�Yfnц׷�<N-I̽�E2�f�R����&�����@	�X©����m��0��b��D���k}G���N��m�La ���'���N1c�W���v�J��-�Ҟ% R���>�LI�kW��}a	I�o��f.*���m��ZY�O'�z[��%e���Jn����vz�H$H��u���"�Oz���-���FRP�=Ht)Iጄu`Q:�����p��ٽ��@�=]��g����-R�N&�ͯА( ���m��&N�޻k�C��ݙ)JK��!j���	�)umx��#X�N���,-�7��.�5��T\���y�	�cO���[�F
+�)J�.�H��'B�n-�Y{��`X+�Xh���0���"�i��"���9��f�0'3Yĳ�&&�XL0OD]ur���޹� [Q����ǱN�t=Q��"#�b՝��E��&Z�1N���"!0m �˕�D��Ji=�Ti*6�z�=ORu�D�Z�O[K!�5�/� ��2��f>��g�Z�i�����l�������2�?�L�ظ��}l�6�/3�1saf��;�OI� �P�E]��g��F~'��|�ϊ�H�%��K9��H`;�"Kb#��V����t��$�E� $գ����upV��R �>���D�Ͱ������m�a���=��u��8Asj����y���!0�{�-�)0�",e�g����_@�|����)�)��`X�ℶ��!8��d6���
�������9eXBqz��޳��	&�y�v���D�c�k�3RZx!�|L�(�x������[��<�D�	ԭ�,��q������KKgmq-QaD�_U`{�M��*U��}��zg��ez�ҡ_5�Ok@��,���'��k ��%�Yj<Bv`a���
'�H�p�y�<␀W]t<�8�&bY�F���Y�1��[%��@�ƙ��>m��FR��K�D��:��C������� �K@�2 <�A]e�6���l>�h*Ht_q�YX׬�m�A�D�z����=���Q�r�(CKd�.�,bH���RB���@����b��q��3�.����P�S�Odg��k3M��<Z@��_01B�k"@<�|H	�e���P�V�.},ZP�0�G��$%�[Bt=:�N�7-%Cґ���'(h/��x�� ������(�bIOXV�"UVʞ$K	j�HV2��R���
RZGVv`q&�PZ@A�ą�LG��+R��G�>���n�o1�-�
A�!'[`M����u�(��v�OP1,�� '��jJF E�-�G��-�2���@bӴ�5`ke$���'VU=�LnRq� �_[}Mm��TIݰh(��P �[�4Ї��l����Z������{m��H�me�:Yq3|�.�
�!�ՐD��R'^��DsrfĚ�f<�q�sIee-��R$!�������'!o��R��^�������1y����'�K��X	[��4CK�B��g���,����)�i'y�ʺ�)@>�z���P��)s��X� ��0�m�L���f�!	D`�6���5��� x�W�=w���c۸�0'�'����XC��-����S,�2��bu�-���0 ���z���h���XKN,&P@��r�SY��t�� �A0�s(4�n�X�sk<��u]c,���D�,5�g�I{F�[-K䂒�	a���čX��u�I�%�a͇�糉G��;���q-a�RJݮe��9���#���xOe}@D�U �l��HX��c5e[�[���B�z�/�(zpW,^<�r���ڼ�;k|⓫IǞ̴�(�/�n�oK쳭*�����1OE:_[8 ! +���"=l��f3�;I�y�L��s$��u���P���M7��h��[`3�_Dk�Ω|�FA�՝�S��r�i����-�i�}hGƬ��0͚����@Y�H�Zֵ�y�C��XC���1/�K��Vڔ��T�B�}�%!myR<$ �2,��Ly;� H��K.}>s!Zx鬡3, J��a�@TS��En"i�	@$X�=O.7Vl޶�>�ܰ 	G��V��%�3�aU�Y��]�	�wk��Y�1I���c���K2T '����0����X����'1�&��b�y��5H�e	#�"����a
�R$5�[��鶸�a�"�a<�X��-���l��`c���C�hY��I�)T��z�w^�l�k��m%��@5�1AH)ᯱ�z���'����X0�BM-�)-e N<�|��3B�F#
&R	��!��L[J��`u���lPlgiٔ�ϼLq|Q�Ĉ(�m*��ź�Zv�
V�JS�S_'�L���GTR>��e�}�#�ل!S7L�{��#̭��:��(j�M�&y��G�<�|�0K("B@��[�!��Rz��K(���תr,� �����ǡ�!^|��i(���HB� j�ٕ��p�,���wM���i�yvNzX�"K��I:)W��[;�}��
д�� @�VTDa�q��.O(V���(�YC1
�-�Z
��[9K���l��s!*��Lw�u��щ�s1jՔ��{a%=	u���		�{K�=���C��:�͢D��� ���`��p���%db��Ϻ�����$(������S�͍��>ZUBݥ	�u@�YՔՂFqm�`	=T�%mD��� �@"0Ǌõ��a�j��b�c��ɹ��&�$�	a�{@���%GVW���z͖�BE�qONp]���L��G4J[�lKvm����Vo7B ŭ1h���c��a0�[�� yƮ�K)�C
>G��������|m��j�+a�/2v��k���Yrذd��g�zwD4H������ƾ��V��[&뷱�h,a�OX'��ȑ<��4`�_q�@��, ��P���km�%#XE�E JG�����|Ė�n�ԇQ�x�K	D��Ҥ������=|Z���Rٚ3V���$�i'XI6q�$�o����z�{*OW�k�!4<[*�A�$��8�
0��<X�)�^��/X�I,�Ŧ�y�CF say��\�y�|�!8�&$H��)i�����+֓�)3eOFx���L5O>��b'�1�ee����%J\N�$9���Y��(�	M�#V!(�+�����e�q��OB�Y #!���[*x&dH{��#2�C��/�e���JI��vyg0���"�
���������|@a�$��k�8��*�X��*��@���s��j��ӭ�(�'���=Ksi(�����@�=J��{����������k#!B�ac�IQ���4|����	IƆ%=h�Xz��0�"Nք��"� Q_T�q1��zb0����<�$�"����O�@�.��ne� y1��|�	�xy��!^��4��kI|$��2!��EYy�1��+�,�
G�M�STm�1y�.��4�A���RE�s��K繜w=(���k�HH�C���Y��n�:�a�!�#��=9���(��B"/��k1�x��A�� ���<��+�P���X��=h�b�
�<FԞVU�i,&+k��ƫ^�|1)H�JB���B�kι"��kL}aHx����ǣ�r�OF *%�	I[���j�6�Ԍ3r�Kz:�f�|B@ *$�f!R`�#ǒ����bl�̰]O/�aĜN����B/�R3��aF�(���LX��83C��1�EU��|VXR�㍞c�Rwi�z�}� U͇���-&.I��(/��֒�$
H�`K	^�hU|��\��%gP������y��}h���K�e�� /�O1����IGů����=9o�F�+'�� �t`z��6��<@��m���X���1P��ٛ�ѡ"B$I��N�P��B B��}J��>"/�ɉ�bD�F,E�D*������dkIS�Є LN���qٗu}*�D!�I6e��{"c],�k��J�$�%ٰ_c!G�FW���(��E�"��Ġ�<B0@��5�7T��3V_*�f���6K�- LR���{���N=lj� �2
����qB�qe�I8��ZI}G�Ue5���hs,�h�pv�ѵ��#�P�ue�/���.c��K2�d���e@2 [;N��1t���L�r��"�����k1��CݟXDM_�c�#5�X�RR&��g!j�l����!'^6��� a�]|��+a�"y��G�1P����a��H���	�uS�⛺��a��<���X���|������Y_l�������&\ZF��P�� Z�Yce'�iiН\HxW��y=	�##^�����2>"'�IOR���դ�K3I^��MZn��NIq���g]s���q�β9$�I-ZK�� li넖��c/�;���1) c%q-�\R�|�%&�C�$A����BTA��Ћ#U�� ��(E����\H��³6ڧ �!<���J3��)HR��O�F�sIfz�X��X��$	����;5|�2>��bC��-b*C�4�R >]�ղ��#!�gV�� Ba�b>|qk�iA#L��ǰ�՘= r�-�� ,:ss'.��a��XX�O}F�U9��SB(�R�DIՒ������ 2�gi6�^1�*�F2s�1%<KB�ǋc1J [i"�}�@*��$$!�BKFR=o##�=OaH�VD�� X�yE�ǂ����`x�K}��O��xb{��҃�$�RW��Y)kG;��:�� �R"C��4!�*F�N����v�c�)_B$⒯�K�+�LDkA=����#TH=�w=���k%��Vsk[�4!�<�k���;����<@�c��^wG��t7�
ňL���<C�!��* ��c�<H�6��±>Հ�`q���і4��1(���)[��(ՁǟX�Y�'W���|֔y�Ա�$�$a^��e̩L]hN�<O]���G�{���Č#Jն0���+Ȟ���Æ�Yf롘@�f<)N7�QV��sc�D�4"Ʒ�HA�CQ���(r����3�������$O�OF|H�Q�B8}A���0R,�mHg��7/�}�X	���g(�-^�!�|e3�b�!X�	"b�Hx D��Y��pL=䥲�gm睒	�*g���H0F��v�Ǉ����� $����[ȪOkĳVLD�M���2�U}[[��,� Ai#)�&5�<� �T�����b!
B1�}��?����/������_y��oW�7���$o��x��_������;�������������dJ������������j<��J���� )ʗ��k�/�?�/������LG� 09�q��e������@�_@ A��I2���OV�?�ؗ���&k��n�rV����&�L�5���j�%�m�rѼQ �*����&u����ęT;��Oc.G�r����f�1k�}AП���<����Kng���$h����w���=���}O?�|~��c����o�} B�
� 5i&���_�0(��)�h9S�#��v���]��V巉�gAD���*uS��bs�	��3�`�42pٺ�w�.t3��,5B0"��7\1�°zb0��ٮ2�;U���|�ΐ�"DY	$W�8��>��7Z�zz?-}���ߎZ1R�;�sl� �1�%U�A��}C��)s�
�*0�~k�� �筽v|@T���SN��v�#�v~`��x���L�z@<\\�	�z_.�N�xo�.,ەj�U�����q<�T�����K�b��l&���~
{F �e�$��PY�Ɖ���f�m�!ĊkvB�DFA)	mǔ���6�J#�<أ�E�g���;y�����=Z(�^�����v��E���˶YѲc9���$⚄a��zl��}so���Z�·vmq6}�R�d�C�X$� o����"	!�Ò`/Qp�+��H>��M�?q��P�{�R",��F���[�t�}d�|m�[�NytIաMS������=~O�4dL1N��˦�p4*8�I�J���A�9L��Ի������,&J��h�Mt�z�=Bx��F�[P�AƇ@E�M3�X�N�oyY�������J�w��b��>�{��H�~'a��,��y(�W)74v�g�nS�O�p{ʻ]BkT���(`F󱗾��S- `�i�a�	�0������J�UE�{����0��򍐑)�.�]��ti��2Uln�Kq"��)��_ˍ���{�v�`��Bڧ��g<H�V�e��Z@{����j�ͅ
�������"�B��jR7��6yn�8�Y�Ib��C Ƭ}o�^S�`��F�5&� ��\�@o��������a�:��N�������ۮri=%�	��_�〻�էt��c>�5�Wv���
2�#�Ā��ߛ���3��å�}�&2"Mj�*9�YQ���:�K��Vɺ3JZ.��io��f�`7B ��{���G�R���rǸ�V�?�*��{�9��ClG��F���zX�Q�wvX�\d�2��*IX����d�1��44)K]���JS���h�~���=�x}�Z�\'7%���c	V�� rB*t�r�FE30g���n�5��U,E��ģ����@T����;}��S��'�0{3Ej ǮN�Tzg|��BW��jУ�D����v�O�3FD��\%�p�8�²�آ}B�v+KP��)'j�wu��gH��"��A����B:CZ=}�y4:f�!�vۡ8^m��Q<�\��8��%��U(HC�ֽ@�3��H������/�!:Ts�YQ���K��.ܚ)ZZ�<=/�D*$9p�Jn*���zx.�3w߇���k'����ܐf����r6�,S���c,��"T�+t�X�chGP%D��=���!���[��N���Ƅ�b�˲[�$Ȇ9r��;\���Q� ��&G."�+�c��!��g2T���P�B�4��Τڱ���YM����c�N�L����H���D���:ܗZm}�8��4p��Rwc1`���	��n�O� Bp�F�=���^��v|��������	��8���6`�(�
�) � �J2����o�~��߫�\>��>�_��z�˟����������<�_���S��  0i�����O���uO�	pO�?�]�X%��.�����p�/��8E׆�[��»��$�����~��M�G��� �P=O�a#��k���w�2�/�0�d������ h��@|�?�kG�P�h2.A(/��6*�]cP���x�p��㣈L7�?�%6L��C�験�~���8aއ �*��M�5�#V%���$9)�� o�l�������<�[�'A�<4���r�`��'Pd�X���T"b�@�5�8��������ͮk�4Џ)��ݽe.ܟS�r��r�X�����c:'b�Xs5�d�%kDf�l��<�ںpRd�,�{�ŞW]_+S����AP��g��W�z.P��$����a9I�z1SJ���v��+! �In+r���0�KX2J���ޓ΀g�a2�u�~�X]\F-��N�At��]Sc�׭9��^�Ol�@�Z��zۨ�����d��,N���͐�ұC�㻹���c��}��c��]C�Y�Ӫ�6�`J ��aX�n ��@�ud�_�4 i�Q|R'�L�T�*�?q�f�/�Al5��ڣϕA�Ю�Iԑm�E�rW,�.�d2|�w�BT�1e�U�]�\�pV�3�j��OP	��`��l(��`��pE0�!m�=�Y9
���or!�G�w'��b�E��x�<Oy��
�ZPf-$]�D��?Y��^ ��]�֍q9%o{c�6�?�P��k'�I}P����a%"RH�j���y`����e0g=UO���*T����J�p�x�'Н� x8����Yr������m��8TQB���%�ԏ. ~�r�g���B-On������:!o��SS�0��RO�D�L��2mt��޷��t��G������
���uǃ�Mm/A������U{6#��A-�T�C��@v0����4ݬo2L�5�5���E5:��Q��-V��W�Q�r��+��T��X�*֜ɨXR��[d-�\�l���uR������/I�z�gQC�hϿ\�䉞���!�(H:�=E����J���_l�-Kk�UƷ�I�PB��5�>���N�!e����Փ�P�����T8`�[ɑ�zJ(`5>r0���d��	�9�]����(&E K'�9O}Wo27T,�*�(B7B�<�K���q@�۽Mʩ�$�<���\�\������N�7!"�:`c�^��
�3ރ��%��IA:���!Z���hG/s�����Е�(��t)�<6�%/������$����f��Xu��4>?�
�J��g����t��	�i5�Jt��k_g�d�΀��"�4ގ����C��	���g���q���H]�����_�~~�e���CpM��R�ObQ�=�T�wQR��[!�wwW��0�羇�'�f,��30vϴ=��A����øPf�9�^,�A�`���`�SlZ�u�g
O)B+���w�9��C���9r�g`����+$g��.�yA��GR�F����Г�Pڻ&v�in��E��ʌf�n%㐪>��4�0!)`���wߔx��w�5�`��4<��uʇ�b߹E�a�a��o�\W��n���m� �fU��Kvۍ#\AlNT�W=���ILB�	aw��H�9��a��bF�|�to�Q�X�6h������Jw@b��g�߹x�N ��ZU���ā�+z�nm�Q��NV��GP�ɬ�S`�����/�Ҥ$��<9��0��\�̯H��x�j �<�=
ӝ�.��Ǳ���p�u*Sb�j��]��h�a�]C��� �pC�(�i���բY&�GYQ���?i�&lwYC�V�X}��1�
D���Ã��8(P���Љ(�E ��J�P���	�q��� KD%Ab�.j﬒+�<�o��}]KlP���a�[�݈��(;5��\	:��ִ�x��jm�j��yn_/@�ۻx�H�2$�>n�8��0DI�Я~,�_ ��e7�f�i,��lΫ�Ik@��W�C���"xC�J$"����{5����8(X��J�� @'ݳm!ā>���n����mY�-lG��{Je���.��&�7l,
�r��O+0q3��ʲU�rX��ӗ	��1����]v�R)|a�
Z��|�vQ��}WݤkaX�����T�L�U�p�mEEWx�y_<CR �?PQs,�X�,/yT����X� 2}��EΔ/2\��p!���22����aD.�1��(�y�4��G�B�콚IK���-W3��p|� \�RRP��TO
͗\	����.B�_�U��QK� ���*'���8� /9����~�o�bܧ6�~~=�x�#]�~/�M��s�� �r  �D_�Oj���
 �J�"� +Î"*���t���6ă� �L�+�#�W�z!�4�
���4*�*�*�D=�߈+�����Ot���_t�����FI�
+��q �PHQ �,(�v��_?On��i>T�hw�2�p*=�˫���(+�	��J��D
(E �V�A�@ �� e_m��� )*� �� "f *̂*�Y��	,��� )�X�%P�`�5��� �@`�.���� ��RQ,�
z.����.?x����֍YQ�_i���}h��cY��"�B�JfD���|�:*�$�oČ�G�����S=)��G����=����*��m-#��8!G�+�l��Y1'��Ʀ�w��M[�m"��Shi�5*��EP�@
QR�2J �EiQ�2 Q�A@
 "e��)J��]B!�A�7�����E6�@m���\��U��2��eZ��J�X|KY|�$r�I�3���l��ǝ~����}��Y��B�Q}�[�Xx��#I=���1�
���+m��RAZ@	���>>�:}}>*��Ǯ�)i
����o�^��;���Ŀu��liF
�����/ψ��?_�E�,c�lhV�ͿT� SO�����Z�u���J��oy�}���|�A�O~)�0�[�ZϏ���6�!i���ӯv��e�3�c��ݥY�z��[����p�'��8a���5|Ͼ�|	�B��-D�O��o���>�����O��{���j�6T�F+<�
�X��Km�lp1�	�#TA�O���~��ݥ-)����T�)��a�o�0�}�}a@	�H�&"@�[5�]p�>��*��!s�I�|z�[G^�I�N��>�a�ı'%�-���m:�� ��m������uf�Y
�@9~$�t���3d&�i��>�%����ϵ�*�����E>l�qc5���8�I)O���ǫ>|'m�3�����{�'�m�K����>$`K��>��7��h��;��iJ��C�a���;���|K����j{u��T��B�|�"BuR˛ �m����f�և��~_K(�bS�Kk,l�_0��V���}��q��+�)��T�{����Z� ��?ky�˘��	>_�'��	��6��Y۷�xOS��o���q���a!���j��%�m<u��l�����!9Yվ��wϞ�t���~΂@!������^����ޱ���֑c�_�	�~=>�,�O�_���e�{�ns�}�N%Ob��P<��ة%<]eʛL������+V|�!�F,OO�;%#�� �FR%$A�&d�o����[&�oia;1���R�Ev�_��e�\b�"D��M~;bXt&���%��b�!��b�u���Mc�f|Ie<Ά6�-%�)�j|it��mN��@��я�ʁ�z���2����S�h8��zdAE�{6�˳�ZgK�U��	P�No�/<���_�������ǹџo'�1Iz�.w͠���RQ[Kl���M�_��ﾽ��K�9�;�>�l`/���L��c������|��v,���B!>���
��Ku���ݾ�i�%ԥc�
�DB���O  <z���t��,�]��Br	@�Y�`��Z� C��e9��oa=���̹����t��)�"ER=1�T�
Ф>^̰z�}~,�螤����@z߆�Fc�(]iħ���v~a�1�2'jY�%=
�v�t�`+l����&���f�*�+�CǊ�jV�|�> ���(�������������NYW�-�@x�tik+AhB_��X�[ڛ�Wx ds�����,�����_T����5>������dp��'��O��u��	�����8��.���'�&12ϣa-��Mka%J�����g��<	�4O}j��>��G��$��i%'׋!��5lU	�i+9�W�I|N,#�D���K!8�ƿ7T���#Đ{��c���41����N�Ĳ��< (!�}o�ue#3a��!}u�'��V�p�&O��jq�%��c>�#�f��;3�CbP�3T!���2�~�s;�P��S�����nfv�{69oq��{�ݼk�S��_�q��u�C9����z��1z+$a�j>���`�cmx-#����,w��!<��Ǽ�C��o�������b��C�a0��|��N��H�
"U$+1�HĀ��dW� �BS�ʥ0JJ����7��ԢD�5IS2�D�(���h���'Ր ��1�|��wXr��f�
0��RWo�ۥ��sR���N�Ё'f`�m��t�	F�0��\��1I�?f]��fE�<F|پ�@υz�?_JI��ԕ��P%��u�) �[,U����O9Ķ��	�̣��vd+��a35���,��ƙ��v숿m遊���<+��8��n�=<k��`zcJD ��B}o�/�j(�m�.'�b�"p� ���m���1� D���f����ba�#i��3_h0��J\�жի!mk��F������bH����+�Y�
x(�ʲ1x~����)���qx�P�S�u�|�%����������/�ͷ�}�)F7�|i������P��Cᐟ>�=Uí<(��a<~i����8��!7?y� �iTc�q��!Q}�B����4��Bd�<0������q0M�*�}�͔���K�
�ǂM�(�>_,"�'��u,���\.�����j��q�q���^��u�mBS��X_��w&m��D�#�h+/�eP�9�1,O��fiH�Vô��O8���@%"����3���}Kz�s;���ƶLH�E	;(�8�׳I� &'���N�jjK��3o��KG8�O�ldQ�B_���-�vj
�a�s/�C���N��6�$����[э�,�����[��}}O\�}�Ӗ$>�P��8����X��G��	�;O���R���Ǿ�G�{��:����h�V(�~�d��5�Y��� &>���o�B� �1���ӃC�����>x���0�@ Q$>wϰ�b�<P%�P�'���S�;��Mi��)Ư��|P����)~����a��)�i��1��{6VD�0�e:��(C�Y%=n�@��{w���$��$I4���	,!锏;��ށU&��&������h�v���b <P����e���G�� b��SyG�)��G�C���P5�7�w�_[ z��*���}xz�z��A��g%��b�B�@�Bt�u�a��U{	^���wCI@P %*� &�x�ӓř�q�Υŗ�3��f�}�T[e��c:�ޱ�`��]o��Wm�������ȭa�`zn�cͱmy���;�{�����1)��[s����p��3�4@w��М�⊊�V�0a%p]����y�k���v�3hq=�[�b�(G-ei �\v�S�d�ѣ����Ǘ>�n�#��Yh<�WWL�)X#���d*R�v	 �`��h)@b�"e$s�P%'dls���*��˘�HdS�ȥ�<��u�f�|q��1��놪Ny�φ�/ ��;y�Ѭ7���8���qݢ�fQ\�q�=3<�77y�EAE[3��@R���#���tpM.�I/(N�,�Nv���Jg]�|{e�	���g��W9y;����g]��^(�f�P�"�"�)v�;�G�A��)y��7���(-�{�|q�lw�{�;TR�T�u��E�Sҳ3���*:�֘�((H�$o4�5�\�1��M�����<�ͺ���;T�S'	�F�#��sv��M��[֘�,'�ȋ��y�<��樌�
\f�-g����l(J��Y��@�Bȋv�j�w\��J
v��Y()�@��) ��]m��v�3��̸�<�����9�h��u�13�d]��!�mo[PD;��D[�\u�*.x�u�M�$�͙
^;�bb���<����E �ﶎ̷��Xj�'�(�r����Ɍ�9��"�Św�2�֯����g$�K1(�@�
��x6�DB`�������(&K1��3WHɪ	|[����U�fc��eu5�:��SQ%٘[N��:���]o�TIz�6����$�)�Z��w�Ϝ�m�d�'��2]��-E^�[x�mrvݘ�Ҍ2�����ŒE��Aka�aFE`�udYj�W�S���(�p�p��x!
QN @M��K�q�\q��I��R��`jF���KO85��
�1�Z��+n�����rZx
�YA�0(��V���ws�&�o&[u�׳����~.հb���"��wۂ��i�dZ�Λ��[�Fo�9� �%]4t�awgqɭz-���!�s}��?�����u�?����x�����}�������?���#�?#����o�?�����֍��Q��?��������A�
t�a����I��E�M~��:�U�[��	\�"��3��,N��C&ʋ�[ֻ���y����Jz3gb�?�D�)������|�<���o�~�ð�$8��D!�PU"DпGB	��aC��ʾ�Ev4�����}	���)��w۲�W���X^m�ٲ��`�Tf	����]GM�Z(���Gf���;l1H��f�t�3ÿ9��b�1�ډ"�u��)�^-�$L����^yfY6��W2�v�!����o���~w�~S�_C����xr���o��?~r�}���U3n����f�>�9���h{���#�|��=��]?� �_�a?�S��7�\��ZۯS��ߠ=��HL������0;�Əd�L��(��$��P�/Ӏ�}=i�m0XW�T����l�n�gG˲pb]�ʃ���5����*�s��M�3��#m���ާ�z�<Y���i�'��=��H	���}���w�C����m�7/����n�[}G=������"Ö:�}0	�w�W��g��ݼAsu�l���(����z�W=�؏>2{��S��Ͷ�3Rk� �$`�YÚ����7.#/F[1�
��Y���J�+I�44%	I�&��h@p���7���8�,��i�ZC$ȼ�O=܋�sN����|U�Թ�V��|7��h�'�=@��U�����@�9`O��{�T��fQ�?�x�{�}6����w5]���9l�����̧Rq����O��v�n��������8�To.�5'��=#�>�[�[�Ѷ��{������i������޿W��X�5���7�U]�o�7#o�7��$ҏ��߬:���v�"�� �@q�@�g}����������K�a��H��h����ҁ?<m������a����~�N�j'�+}-�u�-/QU�����/��┃?֣׌�%բW5rX}O>��oF���@��˨����.5URI��9���"42�@�z�\��j��|7!S>BZݳջ���::w�y�\o@[�Z�m@���|k�dC3v�g���F�۪��zİ�; j'�(q���tg�ڃL�V�P��U�6'V�_z��'��tx1��֊`��Al2O4��2�B	�D�Zf�3k���5 M���qZ��f��x�I�B��˹�!�|�W싍��f����j�O?�|u(ka���st^�lRd��Ȣ�6F�{��{2ؽ�bO�~�z�
�4Ƹ��\#{�'�>�-��rp�`��'Ǩ(g��%����HmD�\�щU�1��zԳ������_q�M��;��mKY
�u��o9ښ{��c���Ԁ�n�_yD�\=(�d^2o2�ޒ�a0��x�9��:���A�:Z&)�ǆ�4^���G�iW��f=>!��u�Y�2�$h�Y���Ulx���F:��|�}���^0O��/�����Ƣ�ӧsD��Nz7�D�G�U�桒7Z��b+��X5$e.�/]hm���p�F�����A��`�oLs�����i�h���l�Q}�gD
� M�bz�%+�h������J�)(M5������S�R��e�7?�s��Z�����7<<��P��'�o���X���<�H��P�"���"t��Kf��#�|�k��G��.X�B��$Q��8y~>�`��Ӆ��b"2��s1R	�a�������e8O�+jk<%hR�
U�k�oo����@+�sj-���6_�)��摵�n|���K���֣}rgܵ�9;�뜶"w1⨡�'J�P�s�� �r+r�֙jJ�/�~m��z���E�M�Y���R�i	C���P�.K���O��M��;r>d�rJ�0Ɠ�=�lc�3׳`8�'���a`�cb�߉#��>�8Pq�ξ���D�0,�R�J*豬>�5Z���~��_�<�b;e_����s�W�&
M�c��~ʐ>Z����$���<xy���{`u��]<��Z ����q���ޏf��o�$�Qe$C
g�~���d������r=*�sYr��h'Tf5=r)�	V��> �D�u��^����q�ᓚd8�}D�:��ׇ�|�co�,�������n�2�P������H��t�=pM�=�M�C��P+e�W��s�����5m�X�mjע�mib�ᝨ��5�FO*?tnP�����j���!���W��
Je����3��y���Έ��ݪ�ٹ���܊�^h��jK�2�Z\�OX7绳�\���En
����m���1�R�\B�|�q��H\Z���*4B�	h�[���2�0H<ia	t�+���^$%{\Z��wo�J�ԣR	��TS����m�fe�l'����E��B���٤��Sn�z�3�����Y��/�����J|(�M. ��f�a��Ǒ�U�<���I ��>}5G��J��3��I|KegA<M֮~1�9q�!4���_ې .^�?NJ���ӽ`���XK�ѕYp��]�hDP �k� 8~2���7���u[xI6D�**Qu>����/�?/�!�Bi�xқ��>݁���쬠��������S�*E���Fu�l0�1��Q�T,�M��8n�j�GA��E)9���M�Ufđ�E�A���eu���{���~&(#����E��@ȻM�NN{�}��]���zr��)T��R���ǔ��X��4�Ne�����ط'z��t�*�շ�x^�0�����'<����4��������J=G/CX��Q-�$K�/��p����N���/?���-�>W��*`�i�^�'�ė�v���|�����ׁ�Л�co�r�d}īCE ��5�B�H���_���_|;�������u���e�#k�M�x���@�����I�f�m�9��;.��K��`y�i������b+k ����4]����vO���V�m�xs.�6�~܈Jzo\�&I�ͭ��^�E1�+IQ��f�=���z�ݢ�3I	Q��kXW��W^���	��#� ��@�ߤkY���샲xɵMנ!��
*�dXTY)W�QA/m�t���c<���8S�u3�mσ^'�B~D}?��~H��BN��D�_�۫&a�i%�^ܷ\Xq��6��#Z:�2;v�54&�-(�9�C@�d����@��2�2PԂ P��(r�ϗ�u�p�����2�,w�>�(��a4s��90�f�ae�͔��|�9p�3��$���;n�$�S.�����m�(�������9!�J^�Bsw�ﵫ�5�ˤ�b�J)㘴�Q@�"%(����c���W^;v������sg��B�Y��rJ�Z�k��s�m��Xm�9�zt,1�J�1E$C3�lB��Z����$��OoME�kFQ3&f#ن	�-]��ḼeZ��H�4T��u�6��+������~���dً���E�o&AIEs|9��-�R�����8�g��&'��8Xt�<,��
3��6�S�n ����&�d���ЧX��.�8�v�o&�3�
"��,<�\ݞj�b��1ջu��X�!�g���ܺ�ݜ��;.�cBg�q�-nz-�ݕ�kfG��P&z�t�dK�I.�������G�?������\B_����4��{J����g?���?��'����F�d���L�{L�����%-���H��~������+�LQE��A�D>c��j?�2fq��&�Tf?5����
���0�B:���n�"���
ƯBL%��Eao%�T�,p(��B5ϻ������"�y�^3�8�Ü`�~6?^��Uw���ߎ=0���bt2s-�� f0����CRU5��i�*e�X?��N��(����~^��$	�:c��?C�)� ��މ���7\ۅ������py4j퐺���.h�BV�Z ��ٻ�=�&U@=$�l'upXdxQ������H�%�Nj@��^�ӛ�h҈��|} n�59�wq���޻k�c���4����R��n��!��Ʈ�S+J��AItA�G.E
H���uf5��w�����ҶTe{�LY5DSP^�5߀7 ,�X������CFi�J��H�� �b�~�15��V1"s�����F$�l��T��zj�Yȸ���`ѥ�(�~���A��<���8�\�CP8Q��p��k�wi���T��"�Ս���=��a��q��ˢK*� ���L��->�k�Du����J�H�IB�q�y�?��j�Pre��h	h��m��ǫ4S bl(�i���#�a`���*;�����߶x��e�rRJ<4�T.s�6�5�-���]k�5��1s[(@h�Eh���F*��"�Uf��u�Nꨐ; $'��*DK�˃�u���-�d��UFE'�"��x�(��*�4��d�rK� ��o{4܀|cuSe`��Y��T0ٚ���6۹�������EF�.�GK�˖$,D͗�N��<����B��~� m{��P��P��0� c���0<�a���*��|:�CV�'��gۘG���vR��ʂ�b[�1b ��Z�D�)��b7S\�fk���g8�9��m��c�2|�ʣ3Ϟ����j��a�����n@th�O��,X@Z�:*v�8Qs���CF�fV�5��L8qD�/��DV�]�!�PQB�*c%I?��"e	&:�� �	"�q|��Z�� U�rœ1��d��zqp~�k{8�L��D0����U��e��^2�`�ze|a��k�i���[�m���pޔ ~#���V�"a�k��+�`*��[����%���V$tH ��g(�tsG�`�Pw��3|P<� Е� ұ��N@� Z����4��%�D-��%�B�͉iD-�+:��X�󽼜��drmc�� �S���-G�i��.L���h �SR(��0��RM��9���e�H@vrcͨZ�� ��5
/ڌ��Q���/H C��c^�2@�594���$5=e�)���A�A�D��y���*p�<'���h��ġw�g��ĵ"sw0�h$)3^;� ��Fg�-���W]'V�0���m�H��x�A[XGg��K�.M �v`�o s�6��3�x65ٰp�q�Z���iG��I�1F3�����1kqA!F��]�L.�t�&��g�3�RJ#+���##$��m"�2x���M�2����55K� �5(D��v����ޝ���RX�)3[$���ǆ��vL(KwHss-bE��vk�n٫5�X��f�#�#ʵ�D�d�J-o�n�.��[�3����2Aq�;u�yu��sw�k��a��!J"-�єFH�͞�FLY����g+5�����E@D� SN�/i�:�ယ�~��v�x�t׆�"���f�6�4v��;F��r�MA��(�v��Y���uݝǋ-UHN3B�95�R=��
o	]��y�zr���x���J-���B3�U��DG��Qgl�)��g%��[�PSJDP�9��]�u^_�.�w���3d&W���䋐XRH��j�2���"�033;�5�J]aA�2+k���2Z��ժ��$�2�7��,�;���2��.=���6�.|��QF���q�����&C�M���D���A�A�L�L�$9ȽaM��f[bdE:ᾍ���Y��)�22)������֠��qw�ʸ#3
�,�3Z�*\�^��!�L��aA��T�%QK�C��I�
C�d%"Y�;�{�u�U�B�R�Cf�,��hY�ЙQ��9�d�TY/=כ˞�aW���aR��(��xK���Hu���{��6��
��p'1�UD��B�P�#�Ij͙j�E�AI�M!�s��*JZ
S#${%�d���LTY�U���'�)��	A��%+H4��Ä/xw�(���� ����+�rG��)���������t维�Q�2Z�(.��A��j���*���L�.���oz�ǵӁ2���	���w�RNAK�P�)i� ̌���g/5�ָu�Q	A绅I��3�h���T�|�B�Ҕ!�������8\�M�(��M�6��:F�j���p�!N�b�J@P(�#�Ӗ���\���Q0%%Ȧ��*�i"J�!���*jB�R������kZuwft��3h�mg�5t�扄O}�u���oG��b*�ε��� d�JIE૦Y�Y%Qf)B�)W$\���N���z�=m�^�:��q�yMg�SFTd`�g�2Ԗ%!�k=U�WO�é�J �#��� w�m�מ�o��}��(���&�Z��p���k(����Y������ȒȮꭂ%�R�d5 �@��ʊ�x�}����=����.��)$b(�IZ�뺲�8�#�v2,2��nx.+��|i1�3�ʁ���2�+�*�����xu���_W^=$���<7@!X�w寃5��=]�ʥnX�UNN�C�h
�{����d�wH��%��P�i�x2JDu-�[`�M�E5��g�Û�upa��o^W=v�6�/m�H�<wl�+|�Tt��%2��p�0��y�2B�*���)���H&��wY��=><�h���@Jku��kRu��fef�h�.3����Xd�fjL��	G��G���i6��PRH4Ѩ��!���}=m������uEgvh�&�
f2$a�Zv�����ed�m%�M-II�����4Tfqde�®�����#J�H�n�a�uׅ�#5�����4Rof��7�p�1��v��XB�l=�w�!�P���Q8ܐ�.-Iݖ�.6A%��Ձ�ez�՞
�F�oek(��Vk+�V�.�=��	�AJ8(�c��ۿ:s�r�%�ݭD��29He��~jB�]y��k-d�`^�ˮe9m���qXG�5�DD;Hgdd]�;G[h6���߿(N2d�=��3x����)؃R��t������5�h]����٭h�����u��T�6���7@gF�����D�
A�{�j�0��
2.���J�j�L���u"vJ&K��"�q��Px�|��#a�aeM8fp���sߕrJ�ܻ+V�ߚ���ܽ��[���-$��9��Y�ƈ��z��4O(2ky2Zb@��!)i���:T�����H;aN��Jjp��N��[ey,���QI�AF�-�kY�s���WS�$
n�W�Ù�fmP��f����1`�3�j�� ���5�x@u���[P�����)E.A�Й��!�9"��)� :�@�1Ҭ�'8�3);'�n:���8q�;z���,\����M�3�
���#�߿WYwk��Z�BNnǳ^O��"�լ��j�mk4Y�諝m���TTUaJ�Y�<C�r�j��t��5Ы���@C��V�;�2x@�'{��Yvxwۿ}���-��V��,�t�f�6˦h�K�v"8��F0�醲�W'�V3�om���^��+�2�ǅ�Z�w�,ێ`Tp�:B.P�ZN0��	5m89@'i)�6�6�N���*n�rN1����o#C��Du�tG�55��M7}�G��0���7|�\u���$��ʺ�%AYf-�rْ{o�5�m&0��xu�����w��ݨ������ vșSN�@��@t�R�o"��w�!�AHw��u��w�8�v`�S�^�'	uF�X�����ek/9rb����Eۙ%U��Mp��G���e�g��Ņ���(3�u�f�^*���6�TRw@u�u�@>	�㊉�Sq�tʹ\�&��^�	�7�tm�d�0��mjS �h6�٤ؒ㶵4�Y�9��}�Βd�Tf�n@��m��/�m�n��0�o�t��٤���Ę�ѽ�wg]g&����j"�瘼`ɥ�1~��4���bN2�e{!;�w�Z�!�p\�|ǃ-U�xmW��W}ؐ�;�{%�4)2i6�ʷ��p�[�v���*7s˙�������w\q-n�ŉ1�Fb��m�1��ݚ1.��[lÎu�����w;f��.�������Z�"��))���I��aE-6�95�^0�.��P�!Ȧ�N�Si)xC�+�v�j�P�2@Sd�\Nأ�G��Af	�p\�8NI��d�I��AI��锝u�G>!�oWigڕ���kݪI߮\X�}�{�k��nr�ݛ��+�A�2
vh)����-�6��ǟ~q�f�]�n4e���2��[o��L��4�*,�x=��|���J��J�XU�*�	�� � R49M��owF@�l�i����a[W�7�7��)3ss���L�[��Z*��[v��i�N2�%:�����B�w�'KM7r��4��o��6df��8�L��݊5������,��]�5m"$��x!2!�P�/G$S� �Gp��0���E�9�R�e�9�¶�Xfj�<���W]��;�q�Y��������m<lb�k�4�:kEp��d�3\��r@�I�5��~� �%�\Lb'�4�n෿9��g���O�o,־^�Ac�n���ms�.��|ɚD#�r���͐��w;�RI�`6D|��E���7���g�e$
��P<�:��mZ�s��=���x�<sk�m|ӭ���+�Q��8��鬍O�l^܃)�V�	xB�#S���L��� �j �s]�Pp�:#+}i '% ?e�����}�u��o�����������m������~��ַ����#?���?��^������MS��?�i��鑙����oKO[�_�O�(���r��?�JC���"��~&�����ۺ�{r�!���"ˍ�yj���>���o�+��3��$��k�r�%NX�o�j��]!�V&;*�>�V/���'�S.H���gֽ'�?��b��LdM�T_�E�&O$c�ݝ� ���1C����{�_��e"#}�D�:�8��;R.C�:����s�[��So��������jFfړx/�a޾�w&�+�}} B0��5bKC�z���2A�2�Jf?��Qј<�]�L��[�Fʬ�����B�����}�Ix��|.2X��w�w,T�z�n��e��S��a��##]��q��>��r�A�
�V�}�[�ʑ{������؜L�F�(vD�<��K�>�K�^��;�H���t��ؿQU�T� 9%Z��.GL>s�t�zpB�+��7V 	H@�ˬn0)[��NR�U* \H��N� L^�:�."�p>J�2}�WW��Lx�J�l�z�y�9rQ�'��xA���n�Z��gL}��~E܃�o��zb@)�&J,�y�t���K/2�c��T-CW���穼B��Zn�Q۶(��[qћ�!\H�6xN�JY6`V��G����S�Ԙ�!ki]�L�L�?0��8X��æ�i�I���O ����0���w'���)<�]A/流�5M�H��>����W�r�8��;�9��q��G|�~��ޣ6/�"i�fގ���<V���#{絪ݰj� g�S<G~Cxy��Θ!s��&�>]+�; ;v�h<W2��r;�D�~R.�,��7 M�d�P��]V��"�2���K)�B�YD��̷OVH0�����Z���X��!�c\0��}$o�����5)T�N��M����[�Zmb%��K}b�(8O🕪�aW�O?<0�����hX��/	R������+�_%�1=}/���e��j�
���"������;*<|G�L�=y��S��$��(ďaZ�2�	6���{����M�6#a�.�j{;y�a�'kֵ�>���h<v��������Q���K�����-�� �z�W���T�J���9WOt��2(O(����ʕ���t�o� �k�].5B�'wQx�;]���J�X�gD���{��r٨ׯ���ϗ.��t�eQ)"�H�G�6��r��6�j�^�]��-���)yy�ڊX�7n���K��>g��폢M�e�ӷE��#�^x�D��|�e�(�ָ��,�{d��to=��6�s�+���,Wh��y��q����kМܭ��f�˲�G�����F�8��}IQ�y���*ydO- �O��=#xF2���L�9<��v._Aw,۩4q��=��������!>7���gi�z�F���_�b\b"��)�;5�\T^4�/4OWC{�!�|{�^������)����ٟ�*�z���Uj���<����*YN���s$"�p<>Im���������/���m�؞1i~-1T�%H��|��ݖ���WVW��#��Ę*S�F޶kz,�T�3Ԩ����+���)w|o���J���NMJ���>m��UTGwγ�,`k�B)��W�|�F��Q<�e�	��sZ�=�&��!�)a���('�*�^���{H����V�\��ԲB�v���!A��'҆��[���>E�HC6��f=��F}]/n2�j~b�����K=;����39Fp��jm�����ΙZ���L�:з�`POe�#�q��~"]̑���9��p04��	A�����2*ܓwYk��y܇O�'y���䁊v��L�II"��1�~;
�,��GT���ېq���E3�����fS)��ZpW"�֕*���<:�&"�$�V�>V�% �����T߳���5$�r��$ݚꔥ��{��j��g�vR��d� �3�
bߚ����eL#�!>H1?�o�={��(�ןUϴ"�C׻�;�������
dr�<uH�����<����ϖ��I;(�.
��a���-�,�ҐY�D��:u�#���_�u.���Na�4=��~�o��R���R��p��]��YX������2=݌JPZ��é�ը:K˹��2���>f�S��!j�f4����a4���r����9f���n�2n�������7�ɩ�9�z'~��Vj�e�_�z�N�Bp�r�ش��s�,�"h$,}k<�|�5Z�z��K2�����q��[:��yb�����0kw�
~s��@�Ur'�qQ�8]N�N�o^t�_����?��W��#�i@������O�:{�����??�׷꠿=�?��O��)����?�����?�rD#�8�!�!^�;��c�@b	=�u��*k�g���WG)b�����*��(�����6i���$��#�əd���9�}��������2$�l��X�@���D" 1D$ʮ���(flvʡ���_��w��P39E�����%h]/�D�D�J�����Q�x";/��p�؅��<��~�Y5�G!rzR��#J.1e�Ȯ�8�a9�*�;��G0�&3/�@
5��H�%p	���Jj�����w&rZ@A���C�ǎ����Ϯ턤'��2@Z�M��X�te�� rmv�\���� �sD:�ְ��Ra\Z&ʻԨ$%pĢ�J�s�j�hn!+�#��`D�1�b%z�!�� �h��C*��7�TZ�uRT���߁�v�����'�@e��#7Ri?FLq$�x ����E�R7���],��0�@h�(1`� S�W'�-����'_���h��9��5�ƨ5���ֹ�f	��r�y��n����8	�R*�
r��qC�+-�U[�ij���\K�0��Y�}�> �� ⾚�O�R���v��!�ݔ���6��G�<�w,;�Q��v��I[ ��yf?c
H�
iɠr	��&���J�&! FQs�Um]b����c! �6 �-�Ҹ�vu�#�@�,��� y-�i�*���,z)���y�]�²�0�/b�X���!�,�I��c�iL3U4�Oi��<�B �ա�rn��ed��I�@fp�����9L��q���}���P�G�u�`PҒ�
�}��MTU�R�H� ������l�M�i��Z���7ǵB9��1�l��z��O=���W�<Z�CG�P�P0aT�-d3Yh�p�M�4�����r�1D�e)x�N%��e���Fk�8�� ����.H��i��ȼ��}��H����^��q�%�)��AI�9����z���[�J n@}W� 3rT��;���̎2E�(L*f�/0f���Q��A dl�KX��U�$���^�کiኖ RZj�DQ��uJ��X��d#�a�S���佩�'8q�b��R���	��]��Ċ\! �� � �ᩤ5d Sq��x!qt�DwZI �$��fD�`4� ��1�\+�Վг��$�8��`�8h�m�l:>"��Ƶ�֕P��DF�j!!���7��|���� +���#��~o}<p�[}6���4��[���Qk"����w`~���U{˹EUJ�p  �d7M��up�Z��p6�&�ं@��iJb�o� u���oӤ	��4$K���K0N 3� 5R�L��C��� 2�8ɐ�l;ɩ�#�C{{V�8B�#���xBG	�5.rU�*���o����>�����?�}o����������1��*����.W��D�������?�����eo���\t�Ɵ�}��'��_����?����T����S������y@����������fP�'ֽ.-�������S+���>��  �1�w�¾я���d�3XC`�);���u�C#F��ƫO�ݧ�����j\H���b�U�ܢ�G�2j��ӝ����y�t��ǡ ��������A��V���@ۗI�m3�{@Lnim��hy4�T=�~��SS��D�UU��,k�wiuF���������~3x�n�.�f\wv�ʢ"u#P����L�$J�%��a\���v��+V�-��[�Ҕydb��i��˚�<� �]��7���Wb��|/��.���x܌Zb�ȏev��R�V�uy������Tkø��S�q{��Q�g�>b�jBKƜ��,N�	= �4�a�g�u����L|;z3���}iӅe�L7
�N^����1n�Wl�}�8g~�"��G�'�n2�Y�_�!~��ו�3���ƿ��Q�����[ה�,��y�e������y3١�-�Q��J�v�l%ƭ)G�r��Ќ����}oٚ-���٫:m��Ʃ�`o�s/M���9��^Z7��,�>�dPr��\Z��bt�j�ǃC�Q��&�������NGœ���\%q�&�#sV=�w=�֫/��.�z�t��E�f���<��������n�P1��3ڄ���۟�RW���y���$g�5�:���u��/Cu1�����#s��.� �p��fl��H=��j+lW.=�F�(gfh�'~���G�ݵ�՘�Fj �$9K�?���
9p���́hc��X<K�'"2$[�k�F�7l�Q\P��A��cp�1^
�"ס�0a������>�-�<��sp��t���Kh�cBC��YQ�䯈�q����ҫ�͖E�֍�'X�ͯrH�J��$p�z>�6ww�+��;��;�5%�{1x:ІM������7�Z�e]�	���4��8�$�yZ�o��O�#��솼Lә��[r�����n��,^�ǒojxi�r�1��'/G��y�׭��S]�\�*hF�:P�Aq�qBU��p�A��ƒ�h��qL9�5=J݃�70���7�h��1��DZ��<�/��+�e��u���4
���όXx׃p��;��AUf-`�",�iI��.�,mɈ*����d್E|E;�,V|ŝ��F��+8����Fœ�(��!mG�)�w ��F����q.��p.�D�o��@!��b��{^��JnA���c�������c�^T<��Z�o�m<����h��(;�E�����O�ϳaw�-v �w4�Q��p������"��&v��0�_ޕ��3�Q
������!����F�YIl�)�#\գ��E�_(_1,��kmf;��؉��I���R��y)G��=��^�WZ�8m>T�5w���,�w̐W��G���ב�f6�yEIF��Ⱥ�i�+�k12����c33�'k�ŤH@n'}�U�P���Y Ĝ��1���:%�BҗE�Ex!N}�
��IKnT�SE�ߥ�gT�@��2�aڒxZ��7�<�)���Sb�9��w��c��Sė�����D/�4��cғ3�:],qv�i���қP.��S�K��S�����Btsx�ѵ.f��鞌�T�7°����IS@´��˾/ńĊ̾�ɛ]jUX�E�/UgWL����V�2��(��	Hb/+�[��8Ɣ�&lk�!���T�������@����l�����p��U��4y��ƿ=��D7��kV�T�o	��@�R�������W�v��������F���id�Ga�J� >�mT��-Rq2s%�K�Irn�lb���{��4FSn=�3�����y7��f��3t�j�\�,���A�K� ���]�,�U�Q��>(�[�<�5�)��QLW>���Q��WA�ZV��ў���nű�Ca���W�P��x�e��R�x3�s����0����;0�SI{��Gr��(nm���vv�J��p������`4>�ׁ;��[aLsN ��?!S�z��?��.S�U~%7�O�\�0�R%^�я�pv#�T�\�}��cʇ�2����mg��L`V*��O��P)�d�[����e�M�u�R�E^ҍ<���u���D��Oir��(����J��h&c��^DէIݤ}֮r�iڡᯟ
�W�I�Z�Η�>l4O%Y�}��hKƶ�"��7Vx�R�i���ߖξF��_@�}}}�  ���8}.���Gʘq H#I�B(�~�<qD	����R7:���d_������/�ɿ2��K]��?�4*3����:g����m�^s��>�o����\c���Ɛ�*�Cϻ��ΊQ�~�	4�?��Pxe���8�@�Np�������LD���c�� @�����ŭ��Z �`��F}L%��qS�+��L��c��Ei�L�daʠ|�B�L��P%D���62�rͫ�EgQ��� �g�f|��K7�CW��
�D�PNu��9L0�(�g���#O��"���Q�E�hY$�4Vq|��m�b� �*��s�lt<'lq1�]��CG���9A4USܑИ��qq��I�
nLd�j��'�4�
	�e�6��HVT�/H3��`H�
$�hĦ�^�I��J�Ww�74�"q��R%JI#��ʆCA��)f,#����uB���0U#b@���QU" w^!���CK͐j��@J���A{�P,)>}��$D�]򖲀��_�2�!��.|j�v� �,_1<nq]6� � ��`q����"�X�?B���P��E_��ާ�Ӧ�?��ƻ.��zHJ�ͺm�r!�@t	#�Bk���7����k��>��,�2���
ɼ��#)��u�qk�@�I������b�XF�8�3%��2:``%g�������B�p(�΁�8f���A��p�F�'��f-4P疋$�F�"F��78D��	쥙&�,��	�!Q�/n�FiP�m@\w�&Fce���QN@��a��=�qĀ����EY1G�1V!G�M�H��^�U��8SO7E������8��.NB�����ᆠV����
e�h8͝����P[#�E�U��Pa�H�BT��=6�Z4�*�<J(&^\�4�m �hlF���-gK�}�q0��0�x$�)%L��4d�(�h����s��r��p��Mɏ
w�Ob�V;�hsWV&�4�^,)�k-`��S�(P��� ���t��G�}�O|}�����{_�ߞ��yF<?���Ha	$8�(A���+�t�� 3_�F�x��'�ax���+tI�B�[q��RӒ]Ş�;���t�?}�{��	gI��������z����g~�q���(�����YgܖF�Z��ͷ�֌�����
���*/�zފ���i�� �5�J�XQZW�
�����GS�ASif��/G@��@ҧ0�4�)�#I� ��";@�P% � ��*4��"d�CP��U2��
���2PR���G�&@�D�D�"�PG!�Dv���B�ʴ���!���Qu(*��^j0� 	�,+����|������p��������������_�|��/�G�t������O� �}��#����?�`���_������V����XW>~���g��/�qd����"xK)E����{��L�iCGw�5�D�A?��EE����\��[a��S��Ϊe
z�(�g˽߱�+�v���{�>��҉Os�N�L���k	��8��,%)�G�W=�
7Hn̟
�����78��������H�,��r�Hڥi�;��֒�����S�����f~��?���&�X�Uf��+O�����u=��7د]_h��&g��ާ��eV�}L�W����>�����  �}  ��u�(%dz�)�Ƚ�4t�;y���)��o@�hk�H:?~�_��4�eB���!%�)��.�џM�Bao�;����5v%��^j���ݥ��gC��&�:}��g2m��j��g��<h�H����l��A�U�����k�6|�[�6�����迊�����1Q�1��Zr�L��ʲ��Ku�z���G��
+����E��jr�j�hUm31�(_~����D��_D�oڹ�W=��̽�S���
����+��w�o{j�{F��z٧�4i�n�F~��:�������h2�gv�m�����}�ӱ�}p��QB=�F���&Z/�|6�JWqԖG7���.�99��>��O㭚�H���i��,�LZ�1'��Kknur�1��
#�8r���9��c�s1����f��0�"��c*��\�+9v�CQ�ڱ�wB���yE��Mާ��&NN�\���g�=w� ���O�	���t���|�2o�O�4V����)�í?�ǚ���dd
.�c��������7R?X_F�ꔡВ;�}d!s���|J|F�ds+[��|{z33�3�{�r�����y����#XG~5dN�Ǘ\zU�#i��A
�B#sΦ	�b�7��:����|'��@���W�=�ƔR�B�oUY�еE��/MH�RX���H�L<5��=�<x"a����Aa��E�.]幋P_��?Yx�������U�w��o���sI%s*�u��n��p�Ͼ$\o�����V����� ӈ�����%F�=�s�=�tz��	�`�Sщ��؍|޹�	&7N�"�������j5>��NM.�j�,s���(�w��bWͭ��������q��^e�����,\ך�/�Vh
�\��;L�BM��ʶ�C�%G1�3^
R"q�Yu�s�+,�����{9 �?�&l5�E�Q�wy�e.�c��Й?D����>8>��ꍯ���i)�+�ozi(j���V��+ROc�v4���%���rn��h����e�{Z<�}�DYL'�{�q��@�Pj���5Ǜ��`U�U��_��#~n�w�T��v���3��G⠋m��KL��}m�|U	�_>��P�������{�ᾱt1SV3Oc4Q�ic?Y|�KK;�:L���UeG��ҕ�݋�6���gDŗ���{%=��$z/+>,~`vx5�Y�؂�]��kK)R� �[��Y�Ѯhϋ�8���
�H��fxVVUNJ �����/����y����؁�r_����i��k�Fw���y����Q���>�f�qVp�{ON'C�1@̆w����Ɵj��n�g֛�������
A�r�0¾sE���כ)n��	<�B5��I�*��t��$�g+���ҩ��r�	ς�-�c������-0Z�I�r��~�/lq����r�|��/�%�ܦW%���r�Zݕi2��T���c�ͪ�PB�o;Ai���h��T.ȇS��򦊤Z���,����OO"�*o1&��jKa��a��bź�[��"8��O*~ʧ��,"�J�Բx�HM�m��)���F��?d�!O����:3��\N��-��e��u��-����:�=-*4���cO���q���F�8'K�_
>$�A�� 0v@�`�[^���M�1�D�u��L�d[��K�d�.�bj�I|��G����0�0�GvM�Y�Z!-tX)��ɽ�Uݤ�SU��4z���Z����OC�2+�������>B�����:�G�X��8s��*H"�Vln4�<�/F$Θc�1|�#�t��"Ư�%�y�8X��2|�Ct%��@+��]Qz���(��ə��`ǆ�Ѭ;�u3�f�C��4��qMw�0�r^��C[���{e���J�#��J3������M��^r��$]rPi�Z��B�ಞ��i���ب���s�Z�Q챗�y~��͎wZv��7K�����brΐ���=<�����{��__�=¡�`�E?���������A�������'��� ��)�
�4���b|�RQ,��&�������Y�N�4<U������������z����vt�ͬM��	�0bo:;� ���횲	��$	��I.�����8���.?�mb�ҿ������J�D�N7S4�#K�?�+C�e�X�����x�=��<�G�o��V�:U��ĥ�:�������<]��o�p�5�'��L���=����Q#���gk���qŞS��)xR ���G�<U�l��M�`@S"]`9Us9k��~/�U^��R�o������$a����^�6��"O �)�]���0P�A��
QTSRD	�#Zʟ$��c�3��j�!��
�&"s���V�8��������6�h��AFp�S�t��%�0X�V�*"��(�o/���?�Q��N6��v��:��Λ�.��t?�#���}1� ��A�BԚ�mUJ༐VYD^=���M�x���5���v褥d_c�q��N�C@)3����x���������?��s�D�.��%7Ɋx�����jץ;}���7�>�?��i=B��퍩/��ʱ�%��|W7�3"��(R��H	��1zѩGmv,��xX�P,���B�N"K�W,����@*�Z���E�E%q`|sտ�N@m��h�-)c(+ ��HZ�Y����?����("�>!��W�˼wm����k���_�ǵ}������Wcm���{Φ˶�[գ�^��f2�)��^ߧ��~G���������B�A	�;Q?M�Z�`�㼂(Rv�P�a����l��H@�N�b�J#�h{�M��B"be����/�=E�9�;�pR� �,;B��d�M�D��>�D�ēVMH�'��֒��-!�^�b+�F�C銒��@i���zE!	�4���ѧ֒ͻ3v��NII��I����� 4������d�-
�Ȱ��*����0�,�������\T#4K���<�������\�^�nﻃ� 888�9�~��WB����l�е����}����(������N�/ �Ϟ��_q���:ڸ�s���|����x�Ǹ_�'Ӽ�!	 ���ֿ�����W��dO�����~���o�W����/������w���~5��}������?���������?��`�¥����D�|�%G������B
�D��q�j���'��%?ʹ�P���w��h�� ��e]���f���BO=ڶ��ĜC��.�4S�F���lMB}]T�;���v��ss��4"�z��M/w�\�zq�H'ܛ۬C�������2��Sf�I�_�}B�s�(!�|=:����'��ܱ�#�ҟ�]��A/��[����x�V�� =	���Z!c����������$�T�l�m�������E�N�q��{����mY�.����|>G�?�>�{�沧�Z�Tݞ<G��{�J�c�t�����v���\����B���F�&��[{fI|;���֮�-#�<����K���Hle�سU��J�3�y,��5���<U����p8�W�[Ȓ���Q���aOST�z�%0ף���������$>7HrQ����mu����6���oC4DLV�&2s�G�ڄǲ�C�L]hjOkѯF����8�җw��+`��G��d�qk;��\�'��V��X!>�涢	�6���*Ǉp6_g�-u	�<z�{�_4�)I4�L{$8��u��'K�}j)��3EH��,��;v�?\�@ٳ&�P�J���K�@^-���@��Zmw�
�+܆|�S��G	����H�G_˔b�n����_Ƃ͘���h7�}i�i�����6��Y]�]�\Ƽ��;O3YhA[|y���o�6=�����+�{�C��<��.g�(���͛o�c�[����瓼~�2���
<Z�>����i7�;��5,�Lĕ�6�S]���+��x�>���b��c��Id�^_��4q�]A/F~���
��Л�zwA^[�|�p����9�2/{��"�x�ԓ3ba��1Ȫ�܁�;�*�2/����u�b�Ȼ}�M�p �:1��dn��V�;��$����o)�?p��2�*�%p$���!ZR��c�1^�.�,���7�q���,	���j��R��!S)��n@D�����_X4�Y���{���3�t;K�z{�G�,���8�����D�3=�?�	��]�	~���P�J�@��f[4*�׃���-�篈��m�{�&<�J�d���}o����>xE��I\��F����{���X!c׆6�;$�~���-ŷ�a'�V�,�(4���H��4�]�jT��ޞ� ��4Hj?��3�Z�(�BK�[�b}p9���b��e��ok��Z)�9m������aǏsP��m�ͯMe�A�}U�c�=�^�|lP�L3��*Gr�����&��������s����6'�h0S;��G�lo��=%�ל緺3�DKym�{sO�fs�����܉ˊ��
�^��|���d�����`�}�k��q�,���/;Ov����{��-���-�-��7�d¡:a�o,����	�K+ �l�)C�.�k��G;�ۍ�; lsH��s�A�>	s�vp�%4��ԝo���m�>���'���r3�Z��ē1E�Y���W`��wSZ���C��)���_�>=���ќ髃��$�/�1����L�S_�r��7�,8��9���¹���ܲX�D��wN��H�k^Z#�Yyr|����y�J����	�gr-)����	��}LmdL��OP�>8��U��$��j�X��wpd=7R"��Q���99^�!o�����m�Th��d�{�%�y�wz�;{�e���9N�һ�������%��j�p���A��"=�d������F�+cQz��~՞|e�a��$�H��ど��>Fk�;Lh�ħ]o=��i~4L��f'4(��B���>6���X�AvLS�����s�XZ�m�{�!_Ԉ����l�w.�H���W�R�� 8���@6���럞�<�F�������YG�5Ҳ�n�g�Q௖��}ϼ˩N����`�+8Y�,1̋���ad��̹VMz���i|g��������8�0֫q��K���)v��1AV��Ɨ|�2�^�V�(�p�@�)��ǥSӊ����GKY�^֋��&�z*�Sr.�ri���̋���ț���V�י%�h��ҙDȓ{�H��8T�.�8�Y���o:.wN4�>��q�Tz
p�y�N��D�K�6�.������4)x����*���<�X*Q�؟���v+�L��׀r�o��fD/���\s(d�:���d�Q%J�op*��M�l/�i,�D��m���O L�2�"�h�x	='�������(��?��x���!<|~���3��1J�ϧ��g���I�OTt������z����������(���~��� �zZ�?�a�@�_�~"�$"~�<_� @�?�� /��j��lֶ����?=��������_ſ���k�$K�9���m�{�������8w��K���~����t��{���ٛ���B֜����"?���g_hmߥ����.�������!����\D��XqǷĞaߙz�N��4�c����g��`p��48T*:娔ɺ	���iF�B@��P�R@%Na�P�"S����h�v K���$q�*�ˁ ��n���2�}�>M$ɑ�N����Y4jX��@��\�43>�4�EN?A�$j��A!��@RO��f� ia��N����k�g��~iB��~�g���Y6�>������~��zk�Gi��au�FUƣ-�C�Ұjd4�T��+�7]���C� ��cM,C�xW^��k�hTY��_�{�����/e�\}��O�����5����'�~��7��G���k1����R:v,�2ܿY0���_~�Awǯ[4���1��4ž?O�M���/
y�|�4\mW�T��Ru��=p(bE,����\EլQ��㚤g�*k?�������=z�ood�;�q
Ty�20�Kuc���~��x�o�?O�����H�V�y�}"�Mk]��.ؤ�JH*���4)$Q�A,��a@u��f��Pp���G
9�N7����;�v�e��klN�ya�t����7��}��J�.������'�2��FmMUP��V�JAj�]1«,�X	,����H�0��ҹk����LD#
�!aʣ%��`5RL1a[�I���](�t��<v� 0�!'Y��\ÈjE�x���9�vkAM4|�^���������w�R��?����|�;C�9�D�e��K�C�HRQ�8ǥJ������	@��*��� ���F(|��>�lՂ~��<��� ��8��m�>?Ay��ŦϜت�8�.	�
��a��)yf����������k�� �o`>��A��k"MQ�� t�8�|܌,�3�tj��6��!U�WuP����ML�`Ol��x�"�v���(��S�E!k37�-��|��U�٩�F���]�G3¹gLWfF[=�� ޮ�8FGS~dً�o���b�gU�g��&Z��«�z�i�'�Yʩv��\�f�����Qtf�z�mg:��a~^4���g:��L�B)@���ocvhu�tT���]G�NG}J�r��w O�S3
C��;���3j�(�nH�=g�>���|�'Q%�w�������H5����]��/6qoɅze�HFk�0���gY�v��3c���?ss:=�tn`�g�Y�z��5;����/ ��ܝ��]����Ե�DM�W\���*�j�t����eQ�w.�
�V�h���N8�R�$���v�^Z�C� y�Lc�<�1r:������4�.��5%�r�؊Q/"i�'E'V��ZU�ٛ�*�k��6�@ۨN:c2\M�!�Hl�!#�nY��/��	J��Ρ �L
V���b��v�+��@ݝ�ؖ�u���`@).�4n��u+�Y=p(��`i�w2�5x3#6WN¨1jc.�0Q�b�Љf��:d��}��1lӎ�Un�y�_;���͛u��/.���F��T7MPx�k8ܱU�������p�H���"QߗL�%���zF^�D��������Z��|��[f�Z-�� #��O�}����_������������o���w����g�n����w�3���}�?p���{��|�?O����/��v1�����]���j�t��?���?ʭ���p�q��G������V�<%@a���l��s1����.��X���!-z\��QCǯ������ػ��!,�+�bny�5��z�*���K탌�v}��j�1n%GlEW��x+SX�G�蚹��Fq�9�&�$]��ZR0qfOtBX�wK���C"^�x��6��UM��!�̜�v�WO���"~�^_��f�ݭQQ�Z�}!��__@��oWK�wx�O�$��g<]��*������9��,*}�g5ϥȯ$j���qY�۾�Q���7ͪx�|����8i���-��Y�%�2�r��M�%3:t2�v��=��b�y��r�$O�X��/쎅0��D�Ȟ�,����n�)sa�Ƞ��n�318�Mg�i�|.D���*"|yL"�kG�.�4����}�+�njP�|���d�G�m.�����O)��/�<�"�29U�wi�BUZʘa���+�,�X�rldf����}
��>�sQb���BR����,u�{X�m�����ل�E��vd��z��^4�X[g���X�˘����wG4�8]\�ϼ�d' ���K�����C�\�5���g���k�tĹݻ�!��j��b^���A���j��]���i]����k�X~�d�cy@�]d��r��4{�Ν[��wM,@�GIO/���YX{'V��<F�L}( ��һϽ�B�����T�o���{3��	�y���3�w4�@���7���7t`�Qm�R|%�Os�Zy]�����v�C�e
��˷͖ttG�㱷(?�trD���M0h�祬yV���	��~���ڏ7��J;������ޮ�7*S�M�Z���|�GV�˖ܾ2�=�	
'h��êo�]���7��}7���{��]��÷�D-��2�ڬa����������Y���I��G�Q�Y����;<��6���|�Ԑ$�į:^!p��A��6&�1]�ga�h�ʡ4���
\����(q���&��� +�s�A�:玪���X����P$	FZ������h�nݥ����7>����Hݴr��4fjd&{\nִT�j����ʹl���������� U��Y9��&�E͔��#�mκ�����FM�wԯ\�7�äd��&4ʭ���m���7�?%��������y�8���[�g�n{�,�!%�"��q�+J�<�H\g����:_�l5�`I7�S��E�A���[���%�dXtf��F�L��U��u�^	��(����>!l��ec$W��{�U�E�g�T�Gj�2�(�2A����d�:��*A�V��pI�X�����q�E~���qn&�����:S�K�{���ox�����|C����^�B{)oUpi)o����f`O`�n��!i'J�&�~�%�t�-�Һ�D�o"�g��0�_���'.��Wn�y��h��|C��&�'^4���U>,�)�B���ڟKS�55�@ߞ� �1��mI!�6N %�5���%mꮵ��ܶ�BK���Îΰ�V�*ے�ݑ���\G���v�gT�#qm"���<�Z����;=Ҽ�<d,lz�ã��1�f)��̙̯����j�衰X��f��%��5�j�.~&�n��Yߜ��������F������gZV����6i&���2��}�� c1���ϝD�Ã=��G�J�^�A��p\��hllaM�a�'�m�'�1�'~���Mk@�d�^�M3Ru��^w÷��I�FR�,׶�'�t�,���4��X�,d�u�?ƝO��u�N[���S@B(��v�hXܖ� ��Vu̩T�N�
u�m�/\ٖd��DQ�7ے��>I_O
�G�$�zx��i�����x�M(��"6���<u��t��5����^}dz��/U�}�Op��5�E5%�"2g�z��s��%�rb�ʜ���DM� W��N��� �[^ך�&����3֙��yd˕��_�<�7c��U$\øX>�h͋G,?����u��ϑ�]��b݊Y���3��V��\2�Ht�����*�yWa\z�V���X-��>B�����d�[�F��M��<�|�?F&0�q�A���K�Ɛ]jBE�aV�&�ɖ���	�R���I'z���%,A*y�cpl�dd��+����k�t��>���~h��{�*��"g���n/r������;����߃;�~���������s�}�}�?��@8
�@�W��N�J	��&'�'/�í���^)��M��S������{���_�=���;S���������kA}�y~��׷~�_���������}�k}���])���c��?o���it�t�HR�h7�����j0�]�S��".��:������ +��Q-����Jס������̑��C�����>��G�}��:#^���O�O���O¿DQ�]�_��A��ȩ�ed܆yٙ�@w$]x�DJj���1T��b���7�x��v 
���0����s��.�Y��YLt�"��\e�����x�~�.�� ����{5oP�����e����W7�Q;f�����:}w����j�۷#���>u����?��~��۞w��~��G�F\v�ohʟMx��x�_ߺ����_�V���'	��I'��2��ӵ����j����S]!�'�|G��mo���'����Q�����]�=��~,�{���{Nx��p�8���5�k�d��(�>���ض:�)M�4�5ɺ�k$��tО�.dDBHn�p�^4` �/��s�;|��)����ۯ{h���/�7�[�ч���Y�L�FgB�#ξ��|��}mo�6=����������}$�?��H��o���:ִ�:�-������B�=��u>�)i?�!�׷���?yKX��c�����~���Xm���B�q���Ϗ�z������^�r��������������H���������ߌ:��V����f�R�j{��<�d��<�1>���+�*2D�2x�>���@ƙ4��N���:{��o~���}6�A��I�  +�_�!W#�'F}��(�Y����xmZ.(�~�G}ƚ�͐.��~K�VG��~�e�*��ʤV�C����?6n��͊�x��i��#4]#*��f��dId�Q\{���79�;�� ��	�.Vю�ע�+���n�̳w���-XrQ\;�zz�Q�P��� /-B��5K�rfr�\eK����Or$P�0z�S��2��d�M�{,�����8:�9��#��aͱ&u[��j�j�31],�͛�8.-�ϡ�&8�]�K{�z�5�T�As�X���"���PV�Z9��]靨�8['�_<��䰻Y�D1�UhWj%ũ���5k�;������3p�AL�kj+S[���Z��R��ܪ���@�I="�.d�M܀6�YRܼ"���nu�/LN��wt.���3R_^Z�՝�-�ά���'�CrIא��ucH
�wy4f�͍���Zb�l�l��vu�p\������<.f)���橔xq��z�W%U�mwL�;�lvxh�f�#ko"��,`��Er�V"�}�B�ʪ̉��ڇ(y�/#�uݝ��sgPr�(��oL�n*�c�����\sn$`�AVñm ��}hPx2�*��/�:	��IF����'xW@<"�T��( >=�����7y�3�')+}����Śvݝ�4+Mt�IZu�z�J�+*�1��uN���tnbU�'s�-^��xw�z�y�a��o%�������w���h#��j[��w�#d�8;ރnf������7�U#�3��[��x���g\\�����s��J0���mkVRv�u��w x�d��=�<G�Dl�dN�*�a�+�3d�7׼�ӿ)����svfLe�٢%�Ϻ]���e�i�����P��{7Qe1�w9�Z��:k�;M�yyx���@9�Q@��#�UC�8�R)�:l��fD�v���Ȭl��B��w��*�$��c�22�fq���ȋ��3�Rz.���+�\y���5n�'Y5�V�˴j]a4���v˖s��wK+�W�&&��rW��W+"��Un��NM�����j��5Fc4��$2ЄT�c���]�<��:*�UW=�ps�=S�YA1K�Nf�w�o�h8���7�?��#�>߇�}��~L���_��s�?��A�R?3�{��g��5����������'���h��[O ?�#�����V���s����������7��~����U����&�?��_��W����ޥ���R�&4e� ���ʖDU:��L�@�����$�j��
8�����
��we���D)�r��:u/�.�s��i��ڡ,`�w�N�Hg��5^�t�>�Nwf��R�H���pj��V
���'Dm�V
�ъ	Hty}�ř��=��C-���Mm�yI ��#�&_}5{�@f��,f���?@ >��]|c3|e�Fi�b�[pC�h{%|�ݹ)fҐ�!e_7RG��X���-?�+��#����n~��6;ԂB�I�򻌊_<�	+(�m'�������Ѓ���B��f��b���[<�X����"���0d��֎�TZO>��Q��������j�kV��̷�7��hT�ԡ���sc2 ���"��<hA"+�ô���,a����s:Z��Z�C���>smqNN�[�B����R���>Ю�6ձ��{��r�YR"�W�;�}�C��n�Z�l��6��n�zs��vyi��@̼��q�w�O]Z�.�����0�7{9��f�K�rY���n�v#}�� <^Pw���D}����2G�Ϸ��ۏy�7�j>�_��2w��ϭ�|��3�\ʝ*��!�u���&�A袶��=H�䒗��x =�*:�w�l�6m\�7��z���A�c�A�5H�_Α�B�Dgz�> K?Y�c֖�'&���g$�>T;���v����	M��/�y�'s39��Yz��d8���j��'�P�\��Q�z�45^ڞ)��˸Q�]�U}5Ը/�Qx� ?���y`-dІ���#}%~*"��|�p��o�9?s�o#b(D����X�����M�ٷ�T,dfo�ް�W.�zbT�S*h:W_mk�q�ڇ�Z"��Fq-Er�Vh���4T>R)&�=m�2��E�W�2q��1�z���g��L�Ěݿ��]o��f\�4[�k��k�zO6�an+�4s���˭�O{"�S������7�q�I�j���޶q�'+ʅ���0]9\OQ<U��G����{	ÁQ-KV����e�¤��ݭD�yAe?=to
	�F8>T�@!J�%�BC��S���~M��4K�&�N�'�.1v2��/O�V��aкA5���h������J��ԑtq$�Q�$�<*��ome�� �y<c���U[ca��s���ʻ8Oc~6�D�6(��sI��^��0S��@����Q1o����B���c�ܨ�&r�R���Hi\���G����e{T�o��$ܘ����D�r{�P0��]�5/$u}�f�ँ�o�'c..�Τ��p��t�Y@!c�4`3��,�-��ȧ�]G���KЕ���nӤZ'd���=f��"jq����^�ّ�Bs+�z���fv��z+����|2%���)�b-,ۤ"����\=ǜ�����L\���{�����Dn'@�}�ߢt�����v�i3*2�e%oTz��>3U����uy[��|l.>�/�n����{�Y"�\c�� $.E�ozI����>LI/Tg��-�N\����c==����Cs�F��|.�y��H�ȹ�}�����qj�In�����M���-t�ǥ4���W/�$��[4J�vi24e�n�es|n8\�x! �R9l�ߔ������e��N�VvVg�<n��\5u�'mbe֜#*�� 5MC4�k}1'�`�"4�x��&�G9%���}���ٞ{�ћoG[�6Qq4EOp?��*�f�SH�*c,����"�%;"�euiF_��=�Ɏ�ViJ��>hmJ"x ң�	�G���L%���:�D���?�������!�;��@���&�T�tF�Ru�ˊ>d�N��"����ޯ����Q�u�VaG�W+l;�+$}B�2����IY�G��Iۿ�w��\g�b������d��W���˻�"�I������̭�K˫����s���y����*H��;mP��{4G_>)�z��0,>�����WB/�}�c��È��&�QC��\h��"~���G��c*.������Y��S#�JW�=�if�l-k���U�*sQ���|��sf���D4K�Q��ڝ�qs�P�Ԭa��1~�������)��$z��3��T��¡	d����og��6�R�S�����|��[�J�U�/6�sȑ{��?�N��퉘ݓ�G�l��8�_ȋ��G.L�.�4Vx��>w���
�tg�u@bC1�gn��9����������~��?d�� ��}߼��|������H��f9����0�⁦Z�Ga{�1���%����F�����-n�k�m)��!�=z��#=;p���Em��r#�~�%�Bt�L'_�Z�2���k��{Ł��K����q<�V{0_�'�D��O�6�j�Qb5��pϵC�T����<}~�}~�Sb��YC��Gͭ�w��4"���k��?���!a��Ͼ��MH�QD��D����5�)tJ�SXu��!"n�ehN|7��ڽ�������ǋ}=�o�%�Е_y��e�׵�ޛK�}&�Q(��)�~0��fHQ]�x���~��. xf�8�ό��U1�|�SHuK��|%"�|FJ�������W����ˮ���������f��Xz�`ޡ�6�3"U���[�l�̮�US�ɡ��s��N"��ߵ��d�g5�8�O�/:ӣ�~%�����K�|׾��_{���v����V�´�GO?^����W����kXE����J��]������g�#-�'�vm�u��'hin�0߭��jS���}��O����̃#B��R��XN�Oz����j:���Z�������-?c�3~�\_Ͱ���u�E!����{��9SG���
3g࿥:�MX�q)nz�����J��}�'���>��}d�f�;t}u��b���#�ܵ3�K"1�m(�/Q�hG��e�^z��x�����jG��}=������$����\������9�s6����vo��3�k,���c�����i�{�|�{�s�kg�ÿk"��6�� ]��o�v�=�_��u~|[f6�wt��4֍��j�9 ��`F$T�@>���K���ߵ�����~CC���?����O�G�~����<�����L��풩߬7������O���e�:3�b���4?��~G��c�~	]���A��)�?~������M�f�1>���)I���?oD��=�^O�x��>�����A�� �+�g2��D��O��_�)�d�~A��Q��:�`����	��,�~?�t�!q2j}���4$�X�!�*��/
�u���3	�-i�v��|���<[;q��2��aq,P��z���?�2���[=�L�W���Af�~`���|m�,"5ڕ;����y���~��������솟j'��b����R�K�R�G�)h�g����]����h���_�"3'�	ɚ�����!\�_�ϖ��Jk�></�~��ˎ���c�2�v�&ƌ&��0���a��!W��kwqn����g롑��SS��|v��V!�q�/	a��H��� H�V����M�~�d�ֆ3�v)bO��$<P}�6��ln:}
Eh����|==��h�U�X��6�E�21���O��|骏%r�p���H<�U��D�+1bNl 7�!},i�ρ� ��US���-��Dʂ���&��B�]r*ac#������s���'7�9�)��T�(9�V1h�j3�Drf-��������	��7��Z�<7�_2�@7WE[3�ʃ�[�< 4�����n��t����:���n�+�c�o�)`��vX���^�uޡ�@�����i7�z<���_\�ޚ��>��}Sj/�w/�7nl�27��<Y�"��U���#slD��'=�a3��-��Q��\-o�C�u�I8G���IE��X)�;�����a�H%ۨ
�zW��*eVm*��Tꮼ�PZ[*�_t��ƭ��'�~j����̌}g�_���8�7�o�ƗJ9���t��ᔹN�D �*�����!Z;H�,�W���%�{��=���R�b�{���gj�_su=��/Uء��k�Mi��}Z+'�Q"t� ��m��,���bY.ܫ�N��
���ע֡y�Å�ְ��Ϥi��������������)���W��,F]��GvB3�i�F���6	[n����_1�n�F�8�'0&�!n��d�FR���<�>�[p��K?*!��x!9ލ�n���q��ˮ�V=g��R��iy]��Ly�� �L���~���4��I+˞����Wm��^����(p/��)�RF>�~N���6aBtڸ�b �^�v��/�V��a��7q�r[̚mI�@��b��(����So�U�SO� " �Ë�-^~?B�S�)+ig�r�G)�Z�G�Q���.{���L��d����r9�`��6�S�I%4���Z<�Ko�����E�V2�%s�,NTS��/�k�>�L�h�p���|Cgq6}ѓv��Rb��ͻ�<��C�>ߢ�3!���7��-�,=���[����l+*&�Ӆn, �PƩ�U�Qѳ����Pu��)Kꃭb�v��<����A���g����e홃�͙�ogP*����x��)>0Q��#d�'�h��~�-��D�G����0�(Q�������D�x(���g�9L\��j����M)����^ҙ��1��[6fF�ܰ���H�� ���d,��|+�?^�<��X�u��46��H���1�-1���`<����h�2v�%�A�s�H���p�����-���+"<,��xi��M��&�W��w��gv]nCq��'2���)hB��Z(�чl�NbOeQHܔN�f�P�u����6�┺	����9=�w��� ��M�,ժuԮ�(����&w��LùZb��=���T����V�9����y�T��
�y�j�'4|��c�N�$���7���QL�,��a�2<{8��8����(ߦ�/%�?Wa_f��e���5����g|\�?L)�vjY�!��� 8�KZ�sx� �%+𞌉P:׵	H�֒��zBeH�ga��O,��*b� ��F �k�@� f��������^�de��E�(�U[�^׊��^�S/��@B\��S��`�&@6�9qۥ%�1�3Y	Mx�pŋ;��(]� �sإ�v���j<��:y�W������l��Ȋ\d�l\�P���XC�},������^����R����;m�P��Uh±������ �Y =��o~�Y����g����}�g����?a�Oۇ������B���|������׷����Ī���������|�p��;U�B��ώ:��m�9���]�J��P,��]v����9�jq�v�5�/g�^�|.��D���O������M�d�h�M]1��QI�Ѷ���S���$��ҭ}���_/�E��6oQ�]k����"�������Ӻbw�ٯ�P���\��?�U8�}�����޽��/W��G[t���j�)�,�qH��~����%�j>;u�[=:{ɋ��I;����������~���E�~���}���h���|�}�q���a*}
ʾ�����9z+�p�z#x�(�,�ǝ�V����ﭙ傩i�D!K�ￏB1�nf�j���ZӞ3��HV���=�ؖ��>{{�w{j#ښ{!Ni߷�{r$ǷV�}T��ۉ�w�(b�ѥ�5��n��(��U�L��H�z}����$��]�wi�vٓOk�J�ڶ���b)f�=i�D�;p�Cί�h�J�����a�P?��lq��M2Z�`u�����E���=�{ӿ](-�i���؟��}K��ju�GKvҴM��d�x���㯏K���������y;��>�$QO��W�0�iѢ���헐�?������Uppo�m�������#���X���_�>��{+d˱��	b��"�G@�d�t�~mv�9b5X��ۜ}�5nE\�0	Θ�Vw*}�P�3���`ӝ��S/OO�����������Q>L81>��k�Dt4rx��^)��յ�wd�v:��*���=��6��9Zx�ע�Yz���OJ�+'��ݱ"��)��7w����JA3����5�^�>tou_	��&�hP��OU����N;�V��!0�\vR��z�"b/i]��M�[�Q�ṹ�'Q5��E����g��9�AJ=�0��{�w��mu�3ԷE+7�7�Y���k;��b�tk�r�&�!��N��}�]�9�b���>���{	Y������6${FaF@�>s`'��p�ꨜ��"j�{L<��w��DG���XT�5T�qW>RY��(���*����Mk�fltt#}��a��=qWE�NW8��A�z��<����T��qQN�ݺ��^$o�J��|sLN�D�p\\OV�a"m��z�sՏ2�]�rz��Gf�����W7�w-��}�0Fx"���t���;f���e���T�u�/WH���+��r�8�E�e��څx9�1us��;5W9�-�Uę��ՑY�N�:�Gj��Y��p���k:��T"�^�o:��-��WpaM�*�'��m���Y�.À�86B�o��:����]Gd3&��z-U#0p�{1ggRD��#\�����"^E�ш��M�)(4�Y����������S��Ŷu�vs�r����g�W\Ma]�Ur\�BIY÷}��u$k�L{;9�By�UՎ�у&7���S{R�ɶ�E\�u��k,�b�vz��:(m�RY�b���̼�J��٫ne
&�wt\��u{�����qVTJ�\�L�v��2�iV��St�:)v�-K�E5���j�U��.l᫁��X��k7i�&'���*7��ȳd�kk��&��*6�a!uï�������������wM���u9Sc�w8�Q�qZ�����Ɋ$������n��-�p�e�N�,��C��˄l֓�e�Swwf���񇸅Wb-��Y��X�K�+��㋼���1O�9�Gd�l��]���s�~��cw�jk+p@`eK^����U\�"���ۥ��m���Tv���yAC��.�N�,n�y��{=��2lv;w{��|ʩ�ɽ۶^)Ɏm�0D��}��� wONc�=����]�m�u:��8Q�o���2�:����82�Q�=��{�-q�1G.{5�
��;*%={b�/�nFВ�[3�.�F:n���p�!8��o'e�F�쫞����"�=��ʀ&�CK��ȥ.�ښ�tp��b&����'cZ�}c��������sT���p� b���Vڰ6;��*.�L������"���э�ؕ��MB ���iͥ[�����mt��b���5e"3���S��k����0��{�d�x��g$ʃ5gY�A�PJ�
�gJ��i�v�&�apOn�Q���!�A�Ȩ��'�RV�c#�QeB�;5�g2^���s6 ����:��Q��Qz��	ݙ�'T���!�b��`u-�5c�Xq1Pr����o�eT\�`���td��cQ��o0Nk�V',�1DƼ����@��V��Ӫ:8`a��j�(�W��*v�zfj��9��
Y"&w-�r��}�$�
s$M��:\AV���ڵ�m`�P۽ֹk�u�2avi����e�E�Q��zy���s��zU_���3[�;şL!�}M�;�o��b�HC�6�VMFl4t�.]-���.s�lN_K�I)����n��۪�x(.�ټl)TX&�e�g�W��^B�U�.U��rcC�'w�犼�x�l�>E�^�f��s;6o�DGfE
ے/9E���#��a�	U�!=	#QW[�śAwf%�WA�����3��,`m��4k�;{{-�P��������������9+`˫+�8���w^_^��m9��#�-�DϹ{�w}�_����8���"�C��2���,��2Ε�+��]HI���j����#/n�� U��bJ[�<���caK\���=�
�z��ٻ��\׀��sz�L��@�h��i��Z�i�a���f݃`S���x:��ӎ�9�<l0ˉ��t�/<Ȼ��Bx�Ur6 v�>ŋhSS���ݗ�&�m��0�n�Tm�qz*�R��.���v�\Z�cj.\,��=W�WώኗS��ΘZ��9�|/���9z,�*g_:شt5<E���`��y�]�����<Ѯ]Gv橅4+N�0�Qv�ݱ{�s�a�u�>�8�ći���H�[�y�J�V�����STN2�	��3Lu��z�ӻ�y5�.*�(��7T�s]vQ�O����O3���ޙ����E��٪�XU�#-�������9���i�,5вɝ�Ͷ�
��1ut��Iu���N��Ŝ(��9�	�"������߹�]�s��A��DK���f��VN\m�oM��)��.YN���IR6���\�W�w\	�i��������nݱ��5_�+r9W�N]Fa7ѕs0�Cd'�N_-�>컹��z����D��c�P�4d�j�f7���8ɉd�����Բ�D%
ިɏ1�$���6��BqP{�[����nۂn����U��F�<�zR�v�������'fiU��Wp|�<b� �Ö�hQqw�vw���LOu��׽ʕ�|u4WB�Ș��8d� Z�o��'H�R/s����e���e�yH�9}Rl�5X�:�A������bf�(��CE{��<Sr�~���ӄ7�G�>��U;�S�U݁��5�c���nq �"�&��lH�����J�[���S�V;��7�2��u��#0��hΓ�un���++uZ�1�}4J}Ω	j�/z:3��w$��1�BB9wV�N�%\US�6���&�)Ì�Tκ��8l`QS����E���v���pC�՚�m��#�nKڶkR٫XN
[9"���������Aw2�FNÆ����D��a諐�����O�;`��:�8�C��(Ӏnzq���-oEz�Ńގ�g�e����������^M�(�1o��9���U���ќ����g����X!+"tX�ژ��F*�������}����W;��5J@������5���f:�+n���z�t����u^�P���t h�{�y��	����*�����)�S�W�1j���[=*n�1X�0���S�T�˄�U]��s&W=����ǐ-lmY]q�U��%�v������2���O��6ʋJ��b���pZ��u�Q���軽����)���2g%G	��r�
r�.�ԥ�ɠVY�J��Ee�Tm��uiא{c%0�6�@@n�5=�3a�qј��`��� #�M�i�ؘ�Ov�ɍ<�/)���ķ�f"�!nj����V��>t:��O�Z��8�ǻ�$t�ꎒ�7Q�����
����&�ɓ*��NU)��/:mI���ŀ`2���]��W�ٝs�`jՇ�7J�v\�z�!�.�)�}�w^OC*��94եN� N�Gy3.���m��Fpg<ɇW;[����!�u��Cu:�]
w�`��
�B-ى:�X7uB�H�l*�n,��9����V^<0����R�] �]빃���JQ�^,(��UY��ڬ�����S㈼ԦM^��9v�[��DJ��F0۱��"^P��T�Rg��8�,k�r6�C�˞��/0-�;�G�9�{���n]���Uܽ��Y<�m��T	�:��ݶѩ��ف�8� �7��v�`P:��uZ*j�Y������7��S�i`Ea�;b�ʬޖKb�����y,]�+�P�H]ӕq�il75�U�G���b3���ɨܓw^�[k�T�|(%��(f�^���;��. ��6�&��;����x�&kZ��yF�+w5�1J|�����Z09М��N���q&��>����u�ա̊�z�k^�̪�X�Zٝ�F�\�=����4L�vUB�t*� ��tW��r/6]�vP9'��ʣ�*�{{k;{z6.c���9JOl(�׌(��9���.�)���f�^,U�ы1�2��U)]�H\�<5�kD_R�ꃃ��H��n3�uZ�7.�����a�s�\�B��Q'(L�<�[z�$��cV�/�BT�<�r�˻2�HS��.vv�j��v��BQ�O`�yܠdwz�Nde�fc�Ѧs}N��R���vK�ڝ���C��)Rz��w�E�.0�:�ʉ:c����;�Ww��e�ĝ[��h��"�����Am9h`(����秂��/dtժK(q�����Gb�M�U���%�wN3��V*��o��'�f��v�j(uLe� �
\Mއ��:'(oo'Mu�m��R�@�_u�N��Ç\�v1>�Vq�w,bn�Xsb5�\*i��hELOU���\���j�.�x�F�WU1��2�R��#,v�FnvUJ��s��h���N�+��pk9�1�Xcob�Ֆ;����}����]��p�3U������[AU��8�`�Oa͠�+uV��U�U�qF����/�_:�Q�\� ��N���t��	���m:|�]G93��̋$�X��]�\
������(�|����j�'����r�k���ȓ�)!T,�⫩fFJ���0@6��7\��9u\���t�)��ݳl�A�\�@P�v3M_��̻h�7��G^�b뎺���S���D�C���Kˉ9����6{-g#1�Ms2�sl���\��WS����q�i�8��:�܇�{kee�OkVl���z�.f�dUd����"�پ�c�Ǝc"E�����j����p�³,p�;:�������B��:3cmB%<�3����#�}7�z��I��gv�f��tQ�ϣ�^��XOGnL�N��<����2�Q�d�����uX�zk�l��T���I�TM�s
ɀ^\�ڍ�;tw:bp#Y��l7�8�]��`�Ӛ�F=��Qņ�e��>-��P��r5���3)e�w��̐�QYWy&�$�(㭄��� `�hÄ��`���+���B�A�m�̜��:1r�q�z7���/�P^�Y����v;#$_e@w{G����6O]U�%�ڒɦ��VUS0GNR��9�wa��ű6 �&��1ua�K&bf���ĳ������+c.�9�y�0�s�w���y�xW����≯�v3v2����2�YK�\�%ndk�Alj���g���6gӳ�F����U$�^�97�f��U�u��_���kr6�_h���2���f:rɓ��h�ʬ�5ճ
3/r��Kȳ�Ƅ��gq�ˡب|8�Q�ӂ�,�6�ђ���'N��˧s�����aF=`	��P�"�]��;��v:�qv
�ԙ�2L�HqZo�΋F鋑(�J��l�28�v��ܽ��-.�F\����GA�*��5<���ܦ�P�	�w�tJ�"�M[�'3)M�U1I�:��}3�/"�gv���+)tږ������36���m�AE�8m�ڄ���w@gI�x�ae��.٫��]�oo��]E0�鼝��<*�����bm$�t�Y�ñA��n�g^VEm�;��e6tLѽ+vN��5V�zb���� ����^9��x���c�pLW�檛�c&�	�'ݵ78��pǺ�춳j����e��+s�.��MS���%X�;�<; �W�Me��#���t뮋�W+:,ΓzY5�S�����m���c:uh<����a�3��=YYZ���1�r{�J��kxod���K�}wK��Fv�Zb�`���ر��Op�Gppk�̼=ܴ�M�݃��s���r^
�]q39�U)Fl�b�ݸ���˄�yd>�s7Fly��T,v"L��g-<n뭪5�ݪ6�R��hT�a訙#Oj�����P����oVݻ�������f�f��roJ�9R�Y,i�Nśث����>҆�єt���~3�ķ]��%��+.�f�����PAO�l�O��u����M�)�^��������Ê�f�cj�Y�� �`�W[���Baoyj�zh)�� �E�"�fxT�=��vM���*���A��Z.{{�{Z���\*��+w\�^�j���a�� {��|y���tX>�C�f�:r]�f�D\�ůR�jaX��y��sY����՜����'h�Ú�g*Tn�Nq�����|�L��l��\�mt
SR�XGL�˷qfh�j&��⫩9�LL�[]F�ގ���i�99U��o2���;Y�ZC�x�j+HN�;�'�.�]�L�D�}vb�NE��n�M��z]WEh�Z�8�(h{9US{;0u��͙��9�����ȕ����@Wd�\��"7���ou˴�=[�wҹe��W�ñܮ:����2�ƍ�]4�"E��w#��Q�괭�s���VԬ���ܒ�Eb����2�6Ҫ�p�tu��1n��ީ�h�4�ّ�Ov�����\�wCn6r�W�V�.Mo<Qˢӝ�ok�ښ�)����R���U��u�譸9���s:�v�\�/wUcc�ߕ3Y�i�����՛�Ƣ�s��j����N��mI�pab���):��r(M��p�=@+��90#f��l�l�U_q�d���q�V�p�g�^�jv�d�o�F*8ug^El��p����̛D��Y��hU��&��/t�S�:���<�a��.�f��s�s7Y�[\����H�0���BPl֠h�}c%E�&71e�Y��a�+�m�o�/��L����h�u5<��tiȽ�������
��驨�����ֺlj�Ll�l����Q�/d��%wv5�Q})C�*�7`�{/*�`��[��oWm�e�k�]��G]��g�*v�rT˃��g�Qא̚�P��]m� �3q|0ا=dj��U�gL0�94��*�%tϚ1�l��Lm[**���Cu#+u<�y�;����:'��;a������T݈��C.r������x�Ybz�zl�p梯�C�
���x���*���c�*P&.lu�M{u���>��=i!&1?y�d^�H�==x���lI˩�Ι�~d#�{kh)j�a��;r|�^���p��SLpǳW�ﹷ�*}��r@fkkn����� O��+�=#���f[˾W����㸸��8�^³��:�9��wM�d��u����3G]u[Qe@���}�&�y7)��Ղ��_�������
����� e�7�)ցo2�3YwTf��U����ϐ�zm�y�*��O��T�n�̃N\��ޭ�ʔ'�b����h����tZ�ӵ��5����`UE�N� �0'E]zg��}=��	|�T�S�k���2�<��D������ ^L��"e�Nn�4:���!��Y�CH�ǈ���93:Zo誡�@z�.;d[��V�KW�py�Kܨ-�toz��ӽ�@����Gh2rNc��*�vɪ[��i��wùÜʶ�po9���BN�͞��Ym����ϼ��s{��ٌc�vND��сY�+�3�]Uy�/N�z =>9����H:�^�77vs�޻y'�)�A
�T8[�{+�Y���N�����ɂ1����u�R�zEH�Ά)s:A�Ѕ`̓Wq8f+&�9�=��%�J ��펣@�3
. �5�梧Q}1.�3J�R]��WGg
��X�$�kg6��Q�v	��Rs����_˯-Z�^@\:r[x�$�3��qO�jΉѐʅJ�S��1���&/*d�������%���ɜ�"(
����^H��2Ś޴Tаq��ɵ����m�V�"s'/O�llX��{X�(�ʽE�[˶�jP�zź��֯/6s��Wr�f�diՕыi�2��[�p����ǼR�i���u����*�'2+7'x�D�6���^� ��:+�D�9ޣ��}靳�>��xP�;y"���)�vN<��fk#6��5' ��nE�ld��,K1� ;s]
���[�6���!b�Z�P��9y�O�衝��u��l(���pҟV���1�^��;��r�cG
����0���63�r���e숒˷=�iRK��-CF��T��]��4�Z�b�[�k���+�>�n;�nT�ɗ111�ʌ�N>:uL�j���y๬�[����Ufl�97�UB���Y;;��-��٬�{��p�g@��w'�:;R��n�iUdΘ�P��!Jf��[���{P��'Ǣ&*��#�.=qs%�õ�t�Y�@ԺgK�4v�|'����	��R�3�M��W�.j�A�ި��R�)�9��f�xX6���ӻ.n*VT������Q1�K}|�+����mBy�t��S3�-�}3]8��;��vZ��[uWc�>�S��[4weO�(��kʦ���5]4�����-�s���s@�v�:<'s�{1�eq�+	�}��v��"�ՐC���x�0�o�k�ג���A�ʬsqQ��P�n��(ݺ��R(u���R�̄�a�[�WS뾘�R�S��6S���2qʡfQ0!��3)V�wn�:I�$D�8C���Ҿͼ�,�y^tU<	e�cj�qq�/(޵*���S�CG�w�4A�Q�\�����Nf6�N�e����[C���2{kLE�)�F����|���֮nN�αN��Jt�٩ٮ�3�ﮝ���#�Ԉ.4һ�`��Uk���3�'�ģ��Z�,�Q��16ww�^��95h�4b�ȁp����=�kuf�uw�}�ʥ��1���3��U֙�z�(��k�kׯ�e�-V��ݸ�!l�A�)kؚE<ˀ��J���3| ;�)�%�#Y��E���"����M3�FwT^�{Sx5D�����$���<���<��҉�ˊ������ЕU3����4xF]mYT�/�wl�8����V.��S�*��wv̳n��xa�-�V�9����y�˸����W+8��[�����Gf����ܧ�������NfZ[�1G����f�����ǫwu�v�l���I�N�[j��e�K��
w)���z�^��R �ns'��:�9�]��.Ƞ���DY$������Pv�|��a����1g�m=
�Qݾ݂z�W$����������jr�֪$�fU�B�6
��2�TT΢�r�7W/{NҖ�]�����hR9��]}j��tr���Cٍ�5*l�e	E]�,�.�����bw[�&d�"� fn-��HN�T\٪�w��sn����eU���S}��1։ͬ��@�<�dH��'#�TMGHD-��8�Ll]P��V�$�X�.6��&&j^V��-`�C��t�vt�������suLr�y��z�9��T�eآ.�}���0�Y��n���ݶsT��7wL��v�NT^[Τx�w�dì���J��V�Wot�]��ONa���B�|r��Ʈ��)	Q3��6^h���ѻ��N���ܱZ1wS�b�l;�:�x�oN䎊��[�sx���(�/]i�U(	�1C���VV�NSSӃ8���Q��Z����ޭY��Szr�Wm�u�ˎ8�1����v^^�<B�:b�d����6%ɬ�$���uT�IQU��j!��Q�'�
)����GhY��S;��4g��Om]\qDm7�j��õ`�r���F�(m܉���!���V�.
�Q�^eIT-����.r�V"������{����1�1�]ܐk�U�s��4ٻ�C5OCV
�������t.�1#z/\�J2�NFA04���c�U�D��}*����7F�q\2^�űz�Dt-������gFA�UpC��ӷxsF���q TM�8qT�X����ܒ6�ik���I�OE��:hH�������5J��VBHX=�Jj�d���{��h��t��y��FfT�İd�>�z�7&H��U�l�=c����]�A�<�%(�&��U�t�������0ž�d���WmdZ�}:!�9|�9��T�F�{�eU��ˑ�*h����3�M9�tV�Fq�M=������	�]S�1mJ��ʞ�Q�/zc���-�Q7Q6kr�l����f����yz�ʋ�71�J�e���fӥ
Y��9�-���ݐ=>�@���w��̱�^\�:8Ν�69[�R<�S���:a�]ٵ���5����ж�k��.�����rV!{}������l��"�X��T V�]�v�ɻ4t�,��@�J"O�*��Q{Z�wj`���sRp|����5�N����W� �>Us�9�&WE��Ci���KOY95F_o^+{�F�;5wGo\9a8qѫ	3;�q���=ф��j;����2uq�UaqQ�b�r�LS7�S#mVi����y�R�x[�6�`�k��G�N�]	�h�{���S����\!��UY�O+�̝Uԉ�����j��urN.�;�4���:R�9p���Gr�	NI���B]�.P�:*�:��#-��|��ܪ�C�'�/m��P���Qj�	F���B��S�z�W'+���o%�Z�gP;f��w.ܻӖa����N�5q#YZ��nD��S�����5[���o"�[��9�X#&&n���Dۉ0+�Sfl�Q�+N㢲��N�A�����ej�ԩ���6��r�e�gpv�u<+�V����RlL���X�b�;�Ӥ��Fv�b֡�y,���5n�^�]j��p��:Q1�j��-�*��Ls�B�p�rp^Vq��X�ɤ�f�#�ؒ �.f�����A�{}w�y���Fչ1C3^db֫��8 �Қ��ּ��z/nTm��[�KN�vKEV�I�9F����,���4��}B��M}�T����F2z4�ufŹT匟m�v���w�wN��<�{Y��}8:Ѻ����{ns��Uz�&�9�L;���~hJ2&��sՙw�]�,Q0�po$J�55=�և3���K�'�US��ir�eJIċ�����U��	���#�)�y��'91c2�c��*�nÓ3x��d��x��姥��P�����&\�3!�z{S�C ��͡Җ�����Z�Ŝ2w�X@	�)�bI�+������F��%���l�9L�ʊ'%L�T�1�&�w�Xh�0Y�n��GU�s�C7;\�j�ӵ
j6Ԯ�d�伬����΍�E1/'�����j�NЭ�Ȋj�^VH���x6-i8r�^��2�ʼ���5b�f�Ctx48a�����*f�3��j╄�B���NgI��Ԋ��m%����ӱ�mrIa��p�.��-"xИ}3 �AF��k2]]]&��{��ޓ��o^�h���T16�s���4\-YEU�±qy+{gh������{}�m��Ӣ��~e�V�+��Wmƫ�e�v��ŋn1u#ye�p��q�o3n�Oer`弽���,ܡ��2�u(�|�ƿ/;]�+��PW�s��ٯ7	پ��9�.pg��tUR֡n�̹�W��Y�m!��EWh��$���&	继�-&c9S�����3��\.FfSu�.^�A�^Wt`^�	�5�x���<�&��ɪ��ūH�Ϣ}�AW8Ƽ�}�{�FT�:�:�k\��0��X�g��f�oc���Xr(fGB/s\��\eP������-��
{]7�o@�D��oyV�l脔��;�wL���:M�\�P}�EU��|^;Uu��nz�5lּ���_J뒬�8���Qn1k����:'fTL�`*P��pq�^��S!���\�5a�~�O��V*�%UŃsrԔսf��bD��2����������t��P�k7E���/W,��Ӽ}�8B���kqZ;j�r�)JVb�3q�f��@������(��'���/h��4�>����`fm/�خΎ��t���kN��.�[W@��`��{��w�{�e��
��{��Wgj��uZ���V;5]^N���E���e�������!O�Qpw�C
��lfҬ3�Kv��)>�V�<*���-���Τ�&
2��v���$���s7̎��� .�y�����{"��M[� T�9�ě�ԑ�Ss]wʼ1V�K��Od�%�����I�5�mT���{K�n���&�.x�a.�Xϙ�fE�e�D��ou\��� �n�1���Pη*g���G����v��\4�I�fC�%��i�ݜ�>�mo��7�e�EF'
����˽�G�Mp��콵��Լ��c�� �d��ռ���ٳj�����5L<���pQ��T7Vk1vm%�M�y8��K�8X��WO]��`WNVͪٛx	��Y�B�31��SmM3#)�TwNg�
������E�`Vc�9�w�9lųW��q35�W��͍�B���ͷ㝷�
�
�$@�5������}�ݛ�Dͬ�+����39��F�t��k�&��.�F���Ċ��f�scV!<�s|��^����Ga��t�;�VrgN�'Ѧ��=���H;)ѤDۭ��G��r>�s�c���8c��W��Ȓ�)4C��]"�KK�Z[p����fI�]F���3��Pm��"/vX�R�F�&e��9��F��3�q�����vK�
jF����F cZ��fk/b�wux����M����E��{��ꦻ�\��qg8������O��'u�����xM
xFk�+h��;<8��۸�䑭8�7ES�vFq��K��v�ZֶCF�C���hɫFa�x�銛'"�w	K�]/�� u^�����
��O=���(2��z���h�����G#+���NLp�#^fLNF�Q��gyɎ��8�;�I�:�F=�S�p��H\mj2Cw�z�l	��H�*��gH��2�6��޸�U�����몓��g^n�0J�nܢnܥX ��Jf����Le�A�h�m�6�A�9+3z�0t���w{]�Wnڒ�S��z�m��JB�5z�BviqF�s��
Wk�7�zM��	#�n�f��t�$am<\sw2�����qu+܋=Z��~^�ݘÍzj���˵EY�Ǚj)G��*4@�ꉾ�G3��>�TA��u�۱U�=R�R�JhkQ�On]m]��ޕF��r�m�Z�Sw<�z��FN����:��K��M��;��hpv�OI����󥙑��"V�.�Ev�S8繩�S��du��㜸���OUp\ڻS�K^���b��;�<������3&mL����,(����"m��K
(�M����C�"*��{2<��J�0�B
`�!��m���a��0�s3Q�q_r}������
���7������? ������������!'��
����%<~����z_�P�ߕ�K�w�I�C���,���������>�D~�4P��}���?o�7���k�=�#��?����X*�!7������  F>a�EVy��q�������O���7sxu/��F�6^��dy�NI�k�g`��:���
$��%���0ˬ�1jk5y��(4�Te@�l��O%�Ϋ�3�tmSU!y����v��&�����EZ�����ڏ��v�S�� _F�Ǌ�!PpO�~�{`|��(��2-�+�E}�ɺ�+>;k���=�+���~/끸U�)-�C1a�W԰��x�	��I��[�]f��/�N�a�9��ʞ��	����$-"	q}�{6�Dk3X�4��۳R��<�L}G�|�1���68��TSAM�e��
٣�O��Ӟ�uq�5�����m�"\qp�K1:ϙ�<m��3�v����9WC[�ʨ��'GQeb��C�>]�"Z𹝒$L�6���45��0̘����I�^���m����Y��Oڲz�u�.ANO�Jx��|�Q���)�����7�3���V������7�	�E~i2\�F(��V<bk��IG�Q�.�H�5�v|�~:ar�N�i>1۰���r9�x���|I����-�e¤r�Z�`T�[���?d�{��v�v>|�buK�1e��>i��wZ���:g��9iwU���"c��;�1k�뗒ՔԆ���"���miȐ��,[��N��/\��|i��^�-b-H�0e���N]l�P���p��w���4&��%�V����)'�؛LTB��"衸c�Y+�쯛ɉa�b�U�l�O�#���\SR����|�sW�ZXp�?2RH��ά�GaQ�ZN��qbB��2����?����(�N���C#_�ƿ0��u��FEՉ�j�_�� �D����#�j�:�I?��/��®�-G��[4��\�������K�6w%�hQ��նbp��&���� ��ک]��{0 OpDs�z�����0eO׽��n��j[K���/�
f���X��t�������#���LFC$�hw>p��a
:Ω5,��a���"�C�v"���Ǐ�"3i>b�5Z�����K���.t��]#�k�bW�5���1ja[f�9���b5:���+�)ph�B�B�C��woL��kT��aޔ��WW��m��Z&Q�����<�2H��zFF^L�E5�*X�k�C�|x���b�-����ux �h�����Rl���t>y����Ev!�=�����m����j��v`�����{�y`5�(�؋��oI�̝��>!��� PY����&b���+~�ҽc_m_{�筂��Ѿ�����s���Z�6���j���Q�{vO:��Q�x�]-�83	r�'U�P(n����2�1����u>�j�&�hew�����`�̉��;r!RnƵK3aH�-�LNΣfj��	2xAX��[�2gI���'o�[�_���O&z��>o2�3��ԲOZ���4�C�U�z�¤}��}�X_Kڲ����ir*+|�;ˁ�v���o@׻�Im�����ڣ	x��d\aW�_���AO��� y��_O��+ f�����u@��Z�����啀8�Ad�4G(s���dg�	7�#��M�΢@e|T��A&^xVx��؂��;�}6�e���#X�G�8�r$�߹N��%�\B�*��q.�F�D[�ޒ�lI9b8�/ϑ���l�3�y�KݟhsF��"��ڂ����jȠ'� �K�fGǑ�=~�	$������*�Ҝq����S��F*�zӊ���q��yu:k��T��BT���`��w&�EW�u�|RܑXډ~��A���3=.E6"��i%�<�n%x(�;��?�rZ�a+ֺѝ@��(�.��5��	�FN��D~~��3��F�(p��z��uaG�5�˶��,�ȅ;�uoC�e�Kh#�)�D_�����y�r��F�WZ[�������i�-���Ǵ�j�X/R����F��2��gQ�ߙR��>w�_~�����k
�"l�*f�	ۏ0�����m�Z��l]�k�{cɄ:��d�sBA
Y+OۻqJ�*:"}�j,Af,�!6��|(������QuƣQ���u���t�CtK�ţ��D��_2،t`]P0e,�.�t�>^5�9����/a��νT�u{Z���EPJyt/ �6𪔔����'��ѯ9�D�e޴9������sTd�Ӝ�56�)i��{��V��%9��L����5�w����.v�
jO۰g'�� �������l_��߯��>�E���g��R��p���_��I���3�$6�0j�Eޑ���zI�z�vU�e�tJ܈��&�������w��eۧ�t�6:�V����S���14�n���M��]�b��ެ��M{�Yz��\ħHԧn�Hvaօ���x|U�D�n���
ZZ%)�GK��	z�6�����Z+S��c�:�4�x���Ǎj�������kW��0U��[x�^t�k߾�6��G�'Zb�0zK	ǋ�׵O�>�7��P$D�!^���J�0�$!��i�'-kE=�����m
*�(��Tڽ���N�x���Uݻw�8�\�m�q�uko/w��� )���ۅ#H���m�Z���W�e�KL!�e'�U�d�ո��u�?i�4H_�Bv�m�RSP��K�+���q��_n����
��ǉD���ښt5Lw�O�5������3Hj��"A���ɳ�B��,��N�</~k�Ջ�8�O��t�Q=���]�9�\���EG ' ��>�pCR��Ǉ-g;��a�j+7�'��o�����'k���?�b@���я4_L9�/���q��k��?u��/�}��-|�-���u�~_�����$~�������T��C�mQI����\}�b9K?y�b]���+��\�M���j_�h���H��G��.}�+�ϽG�IX��,��7���4�~�����~��?��o��P��V,2����*{�Z���_���^|������3���-Z����r���!�a�$���|�&��P�9~�x`o�fy�@��;;�)�ϛ���m�&�k����������ڈK�l�<���YO���3�c��C:�,����A-��}���Ea������V��n�\�><Q;��`�/�Z�/���jW���wv�T��3��3�%Z{�u��DO0h[�5؊���ʮ�LW�Ow��YI�'�}rb�cS[���r����	�/�����)9޻�?��q���r��+��.���tI�>;� �]��g���|u���$%>>{�j�d��^�HuT0�w���#�-2bT�W�	|��HbA�nI��i!����.�)��<~�oˊ]Z�}%Ce,����D���V)Ow�:!f;��Zݡ�/�um�IvQzr��	��Z�T�8��@Q5̪HyRx��ƠVN.m�"�ӻ����A������Ac��RM�*�^��+U��D�m�d<*~csX��2�c&�m�~(Z��ƒ��W��}���N�%]6��[QӁPN��fL�LO��U�_-L'��{����-��Eާ���o�����T�n|t	�2%��� %/9�BK�k�w�e=�WǼ(�R�nY���C�nh�_�6���l��-��	��ʘ����ws���LUI<sJ��*��d|�b֨a�ꃱ�r<�mTE�)x�'�o���5���|�PA	f%���_p�1Fb=�lǛ/a�I�
xPm�Q��|�.�@r�7'��S�VN=~�d;�fF�4 �I����.��l"_���9U"p�_s"!�
H"�Sw��@�Dv�Qf�X�>f��nǷ�u/��ߓn����v���ǚ<�� u���AMF���Z��}C��#�"�#�dTR�q��[2t�E<���z|VLOP}0㍌GM��=XK[o�k,=��!�Os�w��=�<McEk/�v����B�^s��[2�}9v�ֹ�i/q�߄�mL��Y4J0�o
���<ˀ�'p�Ǭ���A��t1Ǥ�c?n�l�&�N��M�L���.q�Tr^�	���b��v�u@�Vۻ��H��E��4�$�Ϝ��cE��4��뀵N\����;	��b�b(�HE��$PX&Åľ��yH�o�)��B�t��x`���W�&���h��yb:"��-��}��Gվ�ȋ5�u�v3/z�w���|�h˽��u��b�P�¸��%���{�)T��a ��;_+��[�= |��V<%yy=.�	�L�YF�s�sJS�<��Kq%��^�q��]�ڭ�ǖ	�z�e�$D��E`^K}����u��
x ��`@�O�}��ԭ'B�J�K�E�z�BHa�Y�Oc)%�\}����%RD
�U{ol�R��q�I���#Y+ZqR��K�֩�}+��J��O�ncw"J�g��4�o��i��z}&�h�4H�`�aĮ	˷-�Y��h�Ω*H#;rz����-�K�0�\8���Ẁc��F��=E��Oo�~p�L�Q��`Z��i=,ǲ4�ZM�'��o���P�����; >��� ��T*��EK^���a�����=�j9���E&ɛ�Ʃ*4�.Cމ~ĳ�29�qt&�(��%!owc��_�s+����4�t/T��E2�M��%~J���7��{�����e5�u��s�U*Õ�`�ٸ��7Gw(����#�%��#2t��D6_t����	O��QI�Ϭ�Z�L�n~� {|���VM�H��|��~��G�u!�d�f2��89~ܤ�4Y�n�/q���6�A9}���
j���Q�\໩��Ui rB�KՏt0|ʝ\F��H�.�F��qZ밗:TA������9�Fu����x�BN&)�����^��4���7Ȧ����D��
�ל=��uZ�>ӗ������VΝ^-�ۚw�᭭C�Q��d���j׳q����h�����
�*�GɃ\���L�k��W?}u�[�����(`ݜ��'��vj?Y��<�4G�9A�aOM���4~\�V���������#L���d �f���w�c���'��-�����~{{������6C��z&�ί��2�˹\�
b���un��潻y[�&y��Q��w�}����a=x�	�?����#���F�=���,��\�:*D�d���UB��Y�������o���qx��z@U2�a�P�6��F���-M�󈦚t�SRæ1A��Vk���(a��aXę��|x�u㞉�̠�g�x�`%
U��:V�p�������i}q��i�-�F�/	��B=:@֭jTB9��TA�H�j�J�|���RTz�M���T�o���n+����s����ݩ�k;QD�	�J>=�zZ);UA�#�J�E6�&æ�f�e�-�E�G����Zf㘵�y��4�]
��u��ϭ)��&�ɪ�B�'�p�k�l��r��7�B�MF�~�1�ҵiTq
�1kIa�D]�e:���o��<���tSl=��3嫰��Jɤy��
�iE�+�43����s9��T�0�"���{��k�6�z�Q�W����v p��;,�|��ˤp�+}�2z���7��FO~��m���1�e[�p�rC��f �T"2T-�ϓ_(��%���0�}'[�{����B����cg�����a�.`����V�ŚMDƚ3�'�@|��b��Ab�=��d��h��F�ڳ�|���VyQTz��F&f;XBi�
�V��RV/�1m�sd�eZ� g:�T��J���2�Y�./��k\�*�$]-��J&j���j�Ѧ���1AF�}��ȘH �iIJ��]�Z&ќ�(�dR����`��BW���@�gH���atv�}M��菁x��$C�">8��ѳ�p	�m5M��0{��I-������*Η�6��AXN�#1�e{�T�i3=��-��� M�$�yO-z���k�����W@g�.���˙���}k�������L1���Ӱ���~%�V>��&"�����j35���"$ ʲ)"���*�,��@�� �|�����^�g�׺��[2-M@<�EI���"�Sj��~_�9R���s�۽��Ew�~F2d���-×1�*��h��( �ş ���$��Z
������|�iY��S�1c;���Dai��������tT�F�zc܌>���_
E�m�)~ s����?���\-��==�;w����pZ���Q8]O��g&l�,�+V8�#��Ѣ ���0��Ͻ�+y�	���4h ���9��n1P�����x��x}g��+�v)0	��W����ۈ���OĞ��O�َ����E8ې�a�J�>�����Nq�]^�?���,҃�^AG0*�R���I6b¨�Z��B�ʢ�|�cs�@&�Kwc��1tj���nm(�[���k��'tr� ��d������D�\�%@��q~;*�Y8��kWOU��3b.��il��|@�;kV�ރx��E�V��xI�m���ב�E�y��wf�H���阢DPI̓	�Y�G���v��'2fnXs;m���Ƴm������QHA�.���JO���>|�I�i��c�!�c�=�U	�~�eu�E��6�Z2t! !>N՛��;��,~�}��w����T�O�Q�@.w� ݀�>���wk��o���%u��X�'(��E%�\�
��e��� �~aYx�d(��Ɍ߄��芃�?3���@�����J���Q�B���U(R���d���VK^�ʪ�s�����&A� ����T1�B��ȡ�XC�7�@ 0�Y�[W�z�h�����%�(B��a ��h�m �.)c&o�UX�JnVū�t��?"5�W���J"�4P�A���Gƫ�夥K�j( mD�%�I�����G:=i0�Đ����db�jמ7�{e�b��v�:��a�y4k������4��&f�������A*U¬X�cUI�`�j ���g����9|z��7 �,�&9+�4�@�����V�9@
�� ��r���	�]QAb�i�H�I>
`��$������C�O�3�@#q�;,�Ā�5� �Iz��~��Y:�hdjQ�"6�ՉP9.A��	�!Knϴ�I�ӊ�n��+�؅"ĭ
1:?+utf4�j
g��Ȅ��@\�tTp����Z�V�c�����P"L`k�.�^+۾�4����Y�O
���O�~O��7�>?�Q�2M�!F*��z�9C��o�گ�����+��FW�B�MY�(`+�����+�(T��$h���US��/��f5�dB	U���� 3 ��ǁ}*�h�>"uL��%J=�_q
�i;
�B)W1a�'H+�\�ȇ؆DS��CߣSq�t�ib���BUnh��Kf6! $fc�B	 �B�0F7�"��[�J0�C
�B��6�՛x/�Q��L�����Z (�l�% ��BaP��(��UfbbB�U�����,�R���qۮ#4Ù���q�#�g����0T(������:%�T+"���xO�$YvD-�Psv6~`�y@�?�|���DB0]��M
L��!?�j��� ��~��J#��)%��Ar�ג�I8���Za6)�s
E����M�]�,��J��3hux
�Bm��#ࢂh\�A$�oV��l�(A�v,	�
\����<�Ȁ��)��Rj�ɚ3���Am��
�T*�U"����t�*�<�����
~���нQ�|�f�}�g[����dWn, �| dz~]�2�

�*`ևf�XC]Qa�  ��S��m�(+����Р5�*�(��Y��&/�U�v�et�I �ֻ^,��3�<EĹ��oK���@^�)��Y���=����ݝ��S�6|�K�i�ڐ(脒1P��d(�����4�I7��0�"���&�Y��I $G�%F�����F�PC��=17�j��(�A&�$�R�J3(ծ׸.j(rB��4~��{��	c��W��&B�F��ȉZV&M����F�DS▙dN�$�pW�d1�!d2���8�')=-kZ�sv���TX0��)Tb���m D��q��=���o���F�P>*���_���g�FT�O)Y�"�P��2Y��x%
�1n]H���	-"��^��R&���
�ȴG�Š�<\<M�&�z}���	���A@�Z7����򓢇�y{!��/xTB�����a�
�����ژ�E(�Y��%1�OxJќ�P���������w昞�����Ԏ>�q��H��y(B��!��[hi%=���S��yM�E[j�,��	i�[�b\)uR�"��	dA6R�GB�P�Wz�	G�dDN��8�1�O~���B]ҥ�0[=�G�@op��ٳ��@��7����,�TQ*<y\�r�H�C�C3�dp��b��P|el���'�m'0rhxY���r=�/��QUB���B��"EK����m1�Z��*��AH�Eœ�8�"/�'�!���c|lpd���U���s�Z�Ɔ�j�AW	v{�"/��� ��4��9u�O2�r�vP��2)OMΠNv(�f.�LHX����'U��S::�䝑�A������m��[���"};C*A���z�0$�T"��#�;��[�zE�X�� �pu����izT1v��Tq�E�� �ِ�8Ί���<����/R�2)2)W��C�Iuĥ��dՙRa�=K:A��
"�nOy�TM� Ncd05!Ƀ@#Kb�:�c�N�@��eeh!����ݙ�a�=Sg�ٽ��0�A�=�Pp�}QȄ��7Z�!tz)�I�uj�=���KS�5��Tk� ��M6*OJ/)�60�_D�!C �h2$5ftΫPJroR�`��M��U�,qd
���
>�!Y��#���L!*��Sv1��(�i�'����o����������೉ւQ�ǷD�������~���5���H`Id^{1]�|hdM����R0�c.�$pv۵t�ɭ��5Tq�(rW�ZI��Z�`����b����%:�ja��a���!� (Q̈$i�(�#�������B�
�d�8�J��M��&��' �L�J���������%�çw�2�>:�kxA��j���e�
���F�vwQ'���<k��4B�K�[F&�%VW��}b6��n�¨�5%fl*u9����%�VE�K{EmJ�d�~�֌o>�i�"Vx%<�еL�@M�>�h�]�H��^�y\�`鐅��QG�O=6��S��[v�BA�N�F�	��("��Gäɖ�"b��"��9Q���ֱ*�6� S��TDL�TVl��G�I++Rv�E@�*ŐuJ�!,���iA(��t���I��V
ɒ�� ��!U$�B�	 �r��p�d!r�t��r$��6�j�*����VZ�%��,�U@�xZ�X+����YNU'e�NNx�V���EȺEDA�$\���ty���(~'.$e/d����*K�� X�Vy�#�?���fK,	��Ԛ�[
�N����UK8��R��f�|t�PM{�Lܜ�l�A�C�)r��G@�p���Ɇ�#�jU��\��օ��	Ԧ���Q�Vj��z�,�"M�H%�0�ˌ��!�h��)x(��T�T8(%��`ղ��8�`pa\����u"�%(�t�D�c�%��8(b�墪R�/�-��<5�Qb��Mn���XܩQ!�mI.�}�ۤ�n���)���ȁ��̤��������J�XM��1�3@�A���!A��U���*� ΋q��|�>v��J�$lu.Z��d���Z(^N�ѴAn>���Ǝ�6#	�`Kh��BY�`�]�݌�2#]DK9ȅ��>���Ag�],�<U�]"��!�^�UEɫ���[���+����8 *�� 'x��y���^�G]h�"�*�!���`�k�:���ƈl��#��!�vk��p\�<G,���kC���f$������vFv�54�d��!�����2�΢����/J�Y5�;�#�Sԅ�UIP�X�Q5�^��XU�q(~�B�rW7xa���}��C=�N5U9���`6��A��>^%��02s.}E�!5(�&d�SY�ח:���5$" S�4���:�BH�Ɯ�&���������;��3�r �і�GQ����f)wE9�%L���pq�M9���2:vn�A=upb�.��;C�+of	�p��]\��ɠ��PE�g�� OmQ�*�0M�oPʌT܄�"�&w�M�W��yk��BN��1P]:Q�bK��E�9KD�J�z�o:b^��F[��#��r ��K�C"��\@آ9ܒ��BF�e�#Չ"t����a$@	B�j����;w�$�s�⋡�ȋ���|FK��z�쪠� !�l\.xElP�3k2��p�vr��G�!k2�j�����%$� ��8����ء؋@5��!.f�ȵVz*�{ԉ�!�� B�RqOv�;:Rv�$x�,H)���	hs���x���%��-l��)�E�ŵ��/,^�6W�7xh����]��SupG�(����ٰ��޳v��9�OMg�DB�B�$B���:Aw��eָ#Sˈ���#1Q�#���]{(��.�!A�=߼�!v��(�t���̥#��F]��B��A��qus�z!����x8�u��6sB����H����Hb�������B�XLM��t���[8�mg�dTP
�@jB���q �������=$$^��-`j�H,��aB]}�\t��󪳂]�YFQ�dG�l j� �&I�y��z!��P�T��;�p���Y�y�xC�&�I!6��U�8���w#�Q�������T��B Up%���B�*P�w�c�@�c�Jn@K���A�u��4��xZV��u�R���������zU�;c6y6��r*##��;-��u���D<V�R����A�ƨ��b6צ���Î�k��&Y\�ВZ��^ $W~���)tʒ�h�Y �^����D�·[��Y� �AY��D��*�XT�y�E]�
9�b���y�t�A Q6N��C �CoKb5��(\C�e*�z��D��<U���� ��\7Y �R�(��V���m�"XAqd�^龦�MC��7 fx[ꭷ���`f��te���Pk3���\@$<Y��i(�?H�x��m�Z�ݨ\v@[c�5U�;�3�J�9BIE����&l��'�댋�mSLT�S	"Ab�iPZ��1_0{�����֙���B,�7�2*�DD|i C:9�]I�@u�f��Y��A�wր��&����A�����[����𔈸&��4}vep�ؽ?�^Dw@��.]4�;$���9sʪ�\��pC��s�$��V�� ހ1����.Q��.�����`^��WG�]�2�@�γ0���	_�tJ^�J0��&��j�B+f|�9��հ�à�r�3�����ڠ�j���ΰB�E�g[��T���_�����U�&��Lih ���M%϶@�~�8��V��(D"2n�Mre�@���)C�ه���C�K�I/ކ�n A �'���hj���Q9�����l<�\K������n�L<
tq@�;��]S�������m�z�$��0BDDd�q��G�6��$i�!Qb]�e�#�������P!��5ֹsΩ �(�,=��GCH�De��`�p�.�s�:�DT�it�F�<��w�PH���r	qj`�8�Ǵ-���QR�{���M8�5��;��.���n핞��rdGj�D�/.C�i��H?�ihjF�G(.Q����-���j��4ٖ����<��$�m4�׮����TU���2���"��6�Bfj�BF-���@&A?A�s��8:Į�}F3G芠7:i���`Iި\�)-`�<@��b�/za���I<џ��8H�L�7�m��=/�t�!�'�2pv�6��
�I:'Ek��u����(�:8��n`A �F&	��G��\��z˶e�Z �97��� ^L�#\��$4$���"䮺(�PK��q(�Y����c�U�A.$�Lب��]�wJ9ҡ!��[�C��N6q�-g�\K���YSWG($�>�tt�"ͬz���/�A������@"%�v{�Iͺ]�v挡�,$S�խ��$�2&)W��D�u#��+�,*\MoG��%�=c�Q���L�doU
I$�8ښDR�n���	m�r�l�mK�0@�d>O�r��[�l8u:H�5�J�(I�n�XqA����K
;5��	p���:o�<��U��$��$�@�T��b)�ڿ�,YQ�j���%RF�$}e��<M �hUPz�:�<����D?��t$��2��AG>EȻ��k{����(� 2g@o'-<�\)۽r�w�H$�� ��Ɠ�:t��@�h�$�EB)ay�"XxQ�b։+'B,�t�T8`+;{������.+�`8��A�utA�7�;�h\�.FJ�̊κ�U��J�v���sH���-G���|������TwT9�ٚh� �Q9Y�r���Ȱ��>�s�/��J
Ol*%�A&!��5�	$�/�s��..&�<��@GB��l�� �&[�+��}ȼ�*�8l���Cjw^����w��f�OB�aB*���:܍|E���E��\��M�r'-W���c���<Q��.����K��_�Y_S�t��z��u�47M�9�a����,�qP�!�$GMzh(I�#� �I6��.YFo1pS2� .;�:\��1���~�K�0	�����i��4���@@ �d�4�4xm40�_؉'LX��	ħT�8Ipzv���IK1 �;H#���`s*$��	 �D�!D4�V�����`I�����r���!��ra��J��R@H.$;:�PԲP�P)T��k�D	��ʻA��W���w5�D�FK�� ��E��W�	�99�@$W��MGFu-�뎖�P���j��K��Y-��;��鶡 �KOU��%�P�]�Ρ2�wA�k'*B�.@�%�K�Ȭ`�ZDg���z)����]s��u.��r`�N��,4�}9� �/j�%ĸh�,7>��,$,O(y���	$��tb���^��^;� ܪj����x.�Y߅�O���v��v[f�����g����}���\��uH�*�	!M�c�]bx�%�ظ�\�+�)t]��x$���ӄ�,YT!�u�=ꃒ�A�&A't��9m�� %��P���B+qR<�`iY:d�A�;�K(�dq.$���������z���]H�� �. �[���<M����۱�rf�l� �EA�FX��t�t\P��L�A�^�_��������� ���`A%ē�]@\m���x3 Fj�p!(m�	�E��MHBA����5Q=3�ӯ.��͎�nԕy(����
<�hY��� <��{���(Q]+�x�h���	 �	��m��q�>HSz���ꂆ��D(!���PE��u��.״��A ��@�0/ J���.�A AX��̓�#��;*$H�p$]TAN=� ޱfդ(�eq�Z�0;cb<gA��Ш]9�4Ś�n}��^WK\\I]�A"��T_(�[��]T�rԡ$s<5fj�d�8Nҷ���Ē��}��?T�e�QL#�]*���T���5��,rbO���=>]�U^)�Rt�8�}Ck���F̜�5RN��D�	ZP�(AG %��襍�K�B!xQ�P	C�J�+$;�\Ak��c�5ꔺAq �� C�+��,��+uގ�H �7!�(�m��d)�!Ԇ!Ē@Bۥ��Ϫ���@g�\�HA��Đ@�YD���F��D� ���0�҅ �k|���q�ƍ��gNej�ţ��}�pd[x���\la�waٝ�Pe
7@��m��<GY���3�PB�(Q�L��%;7c! PI,��P�9'�$���C9E&̘���$��=:�xH�Խ�h��(��O(@��9�JpB��*UEHb��
ƫ��"h��.�o�ir9!�tQ4�
:\fu���K��yr�Ă��'A��*� ��D��^�	��^I$X�i4���P�ĝ�H�ײ�r��:ϪkTD
Y]�8�J#v��B�nuQ�ҩ�D�N(U
%�ʤ�mW�$�u�ѯ���� (UYK��BvQP���z�����v�J�.DF^�@B�pAJ��2�%;EX!D"D*��:!D���\H	�LJ�BGb�SpT��g���lD�vJ��%���]�o$@�@EQ-�m`!�}w�{&�s$���|&!W��3u,�B(��A�P�n�y��s�*G&�v�U�ʠ%�Z,P�jI�6,�	sTT��yyBHr"  !CEָ{�^l�%'�� 7��(�'�Er>�`uFW\2G!B�A" �,��@��r��'�Vu����7W#�CB,�hj� ���vx�h�9V7.��t�*��5
���g�݃�LDP�*DIywB�DVF ���K����%4f�E2*K��zG�n�Rr$S	FC��R*UJ�b�*&�A�
�Jj��%
)��eBU&�w]	��A �D�
Q���)M��~a�3BB9D>�&�2�Tԗ?r*L�=,�(*�Uz�P5�y�Q��B�E��/;�ѕ�3�Ek�:5�M���T��K<�K�#�P���ꃃ��| @����\l�I�T�D,� �E�=�=�\�JP�Ulr�^Hn����3���]����$А�E��
��M���@�iZ��#����5#�#ɣ�
������ �eU�"
� ?J@���䏤�(���EBH!	�8��Q��������L�� ��
?�5�!9��)�r��ȟVJ!K���>{(���)�V��B�&P�W5V(I
8� ��u��&�b�q$/`yq�P|��~	'D�:���0��Dr
�`�j��K��<~۾b�+B�/(��?� P��[/Ft�	!9��4P�}c%�"MAxS!ed(�R��D$�Na�`���\B�tP��M�r��XP��?�_��y�r�ł���D�����l&dd#�B���MJ(�%7E�� J�����>8va��|���
J��ك���l�c�{*<E~��x����O�9��ghK����I�Ĥ�����e�?C�z�m��LJ$#�-w����.9L_��h1%������2�Q^T��XC�	u��=Y��cDA�z����:��PUT�%6g�{)V�XPl��_��sEM�x~t��d�j���{3�36t��q&��d"�H)(��w����EI'{������M��H5E�+��6֬#dU�DZ!(ʂ�0&H�L�i #�_̦���6��LH�*T,=��A��4Lf��%��J�ʁpf�W�!*���ŉDHZ�!
Z��YЇ�O��ǽ�*��K�'�J��3F�����UWܺ �T�EOV/DFB	"ʐW�X� �َ!(3؀����"�*J��(�aH
I� C��
[��	�鴐K׬�d5Sb$�/s+X��!�A]�{+�9DzR�0Te����
W"�;2�@H�C�x�K�*�ETEB���m�]^%�#)�)D�.{��Z��eԵ�Z�D2�c �D�S}7��H�连�,�Er��u,������Y�X�����tJ��A���x��P�|���U��eD��Kۢ(����gJ}�vG�G�F�e!D
���ɐ=�ST|l2�l�'DН́;�,�������񊱫��z�1o�i�t���X/�Ƞ��$Vg"�p�O&�QZ&�Y����Rl�V\)U;�!�����[+��wk=!�*&U�St�d��3�뗮����,��+�`�@1Q4(g�����F�5W���GA$����u�J��C�e��7k��h鬀�����*���7�J�
(C|XZo d�[b�F{h�*H��$��JZ�r��zz����6��!���$`��E���b�g�=�0�!�5\`�ERȪB�~��$��6Dn'�|�X?����Iv�kzZ��"��D�$�*�"Ly�E��.�5�QxK��)�~M�Y�> ������oV��,(��?2�3 �6���&�.�~��c�nMK�3�7L�1����A4��i)"����| h�'\��g�M����`*�g��n{܉e�2���kQ��{�Rׄ۶@~k��G��b-�'�����A@~g�i���P���u�W�d��e3��<�<3�"�t��0f��AZ>!&dXY���Hb1�J�ug"7aB_n�<sc�n~�
KǄ@�#g{h�UTe�! �C�F}%%(zY�W
����Ő� ���P8ŦE��`*����FX� �_�'=/�%!�}%f'��i��0b�Qj��{��G��Y�F9z��WD/bL   �,*)X2�+�#��;#�K��R�3@}3B`�D����i����}�[�Ժ�`��fC���R�a�o�)t���H���K�+XX4��\�I���S��K��U	�l[(���0�����tH2��,�����8~U�{h�5���P�BY�ʶ��A��@*�p��K�#S�'��Q	҇-edAw���	�.L�Ee�?0�>�O(��E%�������lQ�RW�f%�ԓ�Ә=����*(e�]�A�S���eĉ��5�����Ҁt1�$dPH�����%i:F�̨�d��f��b��'��ya� �TD�t���C�� �����1LPQ�`����!����m�d�_Ľ5+�mX�I8�Q�����"�U[�$?-,�PV��Ш��J�U�t�;¬!1_�s�j���%f���5�L�������Dv�<k3�X� R뇲���ۤtcl'vGg�^T`�r���u�
!=S&ȆG�lY��¢��5W�zl����]]�q��y��T�!&��/	:�Y�"h��:[Q��Af�����1�M4
l�d:a쌊^����[��F�7�2��(�0+�� �,�:6��Qu�X�飂a�$����\����3;����E��G"Qv��y��L�&� i|�!�/~JQ�!8z���a�oȥ"�%�t]2`�FNSU�7�Tي���dG)�"(�B#0��:o�^�2������LF�H:��M@�A7Q'_1ftH� fJ���1��t���E�J&.����%��`S�f%�T�m��s,�i��tP2A0/���5�>G�&�4� �J�)d(7�p��]%[�!�;Z��!"��n������<H���k���(�'(�������7綕���L3�ٛ�I��x%I�2�Ah燷)R�$��(c��we���튌s�N��&�WMB̐ ��/��W<uT�}�ԥ�����;E�@��N�z���WG��$E�P�Eq%V�UxTF��]GLO[�V���S�����������Y^���td�Br2$.��7�h����ob��v	.��-=��Q-Q#-uX��-�ʌ]�we�{#�-v�2��@C�*�3�5��uDD��:DA
e^�A�i|�JUK�tQ��!L��/�ԣ�k%��mT0]��q�P�w��"MaxX��v�B��r�U����?33�k
���]��Yq�]1�B�Ø>R��<�GV⦇��A��8��P�v���)-��rj+j�S2�7��Z>��(H�)PJP)&|�LZ,�"%,�u�hA��h=ʉ�CAZ�(�3ӛ�\��TW�����"O�ħ����q�%�0��֡��
]�*a"��D�5��^�H��w˳rG%9��{\iT4r��"h�"��n^j��}%ob���#��
�Rw��	_C`E,4�L�]�Y)��o$t
�́���By�*m�Q���h�=��]�Ʒ&�b�]2�-��wB ��(��h+��%��BY
nA���*��-"g�"���t8tUΥ1|�t���'%[���U��-@���&���{�52)��zX<� (�������X*%�.��5�=�N�����`J�*@[�%�B���c}.�%�T`.{qN4�d\�wa�p#�
Mp:I�Y����M#����0.m�s�*��T���u��2�_�&�+�F�u�q@����l�I��LM���CP����1���KV�+Z+��*��C&�3fD%*�b�,됗�jHx Y�؈b�DHE�o7T�I~ƴ���L��8}Ŕ��/|�H����/g���lB��S�#˴r��S�:Ghc5@kH�$�FX���:Ժ�c�H\nE0Rd8����8'�q]�>��LHE2I �p�j��F;�$�$��$���7�i�p��&�gX��^�dM�H�.D�#�a1 ��@���ET{�r��+oL`�֥Q���y|�K�j��=�z �{F���ƻA�@��I>8�#Ǿ��;h�hEkt�:a�M��5P�͗��A�快`���l������4�$�'6����B��8�;�Y��� ��&Jԇ+ [�
*K\�e��^��b�D.;&�f����4K�R2��!=��q�$i(����G}"8�`2R�S�	/Lh��Aq<��N;����*r{�%������ _w�G
.�ք 5w�qz��*��fI��䅄JL1��d�:f�`�(Ϙ�����菛��>q��F�x�`�}1�*��Q9�g��Aɒ��.Q	E�r"_�\l�Mm]AD��ٟ���_[j(6�U�/��&]y2�I ��"I6��{�����5�蠑Ђ�[��Cjڍ�^���j�i��k���E�Ut�$��*HΆ+EBF����m0��0��"'pΚJ�%T�u�@\H�ŲPY�@Ahω��0����|�,�����r�}���J����ƘÌm$�FjN�
���n�k��;.�q9�Bf�G�"����#��1�\��N��#����o����閦�E��}
������ر�汶��6����PF"�6z��3���I��[%��HY������ĢW��0B1��-L`��	)��n!Y�W��� ܇�e����k^_L,�\F&�h))f�w��բ���֜|� �DjB�Qӏ6�1IG�x/�����0Y��Y����յV �H�Q��	�a��x/��:\�l�,	���q"M�1!���TM3}�`�0H,��S�V��K���.t��=
q����I�1���i
����,ʷ�	z�;bDl)	�sE�#L�T�X7��l�I��u�Mk���*3q��H�k���/���;>(��:/׿l����\H�[�T T������ҡ��d��e2ƉF�rLza`QR�˙��Z^�KN�J��)adУ��R�A1>� ·l����$�9MB.@!�����2����J�" -D�#P�khg�]��� ��l�E\������ ���&j���B��"p��*�.����"�ֶZ�gܒC�(�|��J�Ērinzw������t������]�F*AE��h�Za����jw�m��`���Ѐ��8�*$��e�J�&$�����r�,�S�Cv\�R%哛�,Q��!	)�&bK�$���8¶�]u~*�XEd���&��J*&K˙H�I"n�X��u�v�w6B�$A�"'��'#p�5�����*�*��Y���B���Ead1t��~����^�Qn�{gZ�h]y��h�0��5}6�X�Ek@�H&�)�)D��[�v �.:t��2Dq�d�\A6�2��P�:N��EK�!��\5�d�0Ґl#�M!k@�F��eG��%^_�!�QBG��k�}Ѧ���;�^rླྀ���5��Fׄ�$�'��@�I�$�yш4҄�Vr *�h��n�GQ�n���]	�$Dx/y��2D�/���TFz*5���}_p�b��ߎ����$��J��Ql2I�W���i�&���3�oPƁ%Ēb�2�Єm�`\�ҿ�$������pWm���d�����=��!qS�� $K_��\��msFʞ0�<-20L=��q��!S��bi>ë��8Iܒ�3�� �#��\�7��g6�a_nֶ|=w{��o��:dҺa��@����!$��=��q5��{>�K�lf�C��� ǭ�m>eL�@$\���ȑ �h�h�ŷ=8ӧ���)��ܥ�m�P��N�̦<�u� ��%�DwQn[��F0�:�M��$�]j��� ���Ѝp��{�:�쓚)q�s�H��:t�xAb8�q���r6ӓK�aT��`��JiM'�r*Mk-4�a�ru�@�'y`I8]8z闾�7T$X��PH&�]��d)a�o����Nn�ɹ�M�⺦�?h�h��uwT<�������yZ��}T���Z��)�T�������@�%v����[�9��ǙQ�jQ�(Ltr]B��z�ˎt�4Dq _,)W ��vΏh �� ��`)�BIxN]E�,G�cG	��7J�vz@�T�5��b��x�>UH���8�IwDM��\�|Ϙ���t�q�ev$ءq�%Ə�����鑊���mP�	'�R� �r��Թ@I(E�b1Wn@.�CqڳQc�[���(�Au���aB�a�Xظ�ݼ��<#���\A'ZeT�oS˪w
�p$A^�ќ'q�Ιp$��P�@'C|xWHlS=�� ���ҹ��+�E1^6MH��˞�"a	q��4��q;aF"�+f��B�(�H:��a�F5���%��zX�N���׿�!�a�1!�A$�4@��,l����!�$�m0���f�t��n�(��W#6�$�� %�j4[w!�}�f"vp�N�_G8��A$���B>�%�
��.G�Q�#�$DM.夬�_��#K���L��w! ���x���7T� �\�� �J�j��^Ո _U��V!�H�`MUrI/�� �g���@�ݩ���ޮ{�(. ��F�?�b6Vl��Δ��(H'<��$�w���<vD�A臊�U�E��H;m���J�tLB"��?R���K,}r���4@K��Ԃ\�A9���8f���(򲻻Jn�C�'B:Q	|[�����b7��c� B�rjA��kD��q��n	&]4������ St���(L�"�$ ����A@A[�� =ۥ��`��͂WnW�t�(�C�-հcΆ|a��k$�r*j,=����1���u���#��$�\$U�׫�������2		 �a �-�9!L�^�(�]pO�= uA&�P	5�W���"� ��C�x�t�<���̀�(b��S���K����<�z�`"\I.#��6����+jZdgFr#� ĒH$���r,���s��� $2��.C3|]���� ��cR�P�giy� �쵃���@qn�yCe$�5t�nFp��yq�Ƞ���G��V�(�����Z��h��"���U�R����ǚ`8��	$u����  p
]I�a#��sH�� �P��5��qN��ͅ�DyOt�SO>Z��x��ϸDSL".U�(f�YH��gU-)��@%�̔�)9� I1E"�� �BI�,���D	�B���E��ҡ����l�I�M�$�R���՜��܉�X���ɐ�~`rxo��7�\˷28�O
�m\��k@��3B�2H L��9��=R�Q1R��b$\�H�TU#j���J��NM�%�|����pA&�Q���l�u!u@�MQ"�EJeG����D�P��^h��A����� �j�
~�+�P9�xj8L���;��Oof����'�����;6��xDs�	$�K�P8��l	#7�h4�8�T�?B��
�R�j�H:����y ��#�&`���=�K�=�I%�5!Gi�,��d��#��A �\M("D�X����r %I�^a�|�@�$�uPT�8AK��+2��8�xn���@B�n=s����x�x�:&n�+�h�X��� A��D *�~��` T$I�|�b@�۷�
�R�<�4� �M0�0xQ�A	9K*�PC�၊���I��΁��?�IDB0�dbH����x��UQ�W�R=Q`E!k�.�+�2�E<�*d�D �����[~��	��oV��
�6D�"(�B���� d��Qi��+�A\\�@x�4�;@`ض"�t���
&(���ʥ�!��4,�
�.ĉ��USG�����7ww�R�uJ 0*B����UM�Q�I�)cW����s�a�*.E���Y�,�l�Dq(��苕�8"!C���I
I���\y &g�.sˮ�Qԓcrt� ���$��O�I\�P�O|�/�u&��JC�$��,ѹ,%4.�!���d�X�R}Q��k"��T� @�Drd/����؀�}ʡUA
3�J3��!C�p���@SeY@��L=V�H�"�-d�RQ�.�E�`�2�8�v����$�K�Ȁ��q�G��>d��4��It�	�!�D薳�A=�-�#�g$�z��B���FB.��l�,�T^nru��p4"�on_7�9�33���aͳ�܇�hƭ��k�zI�}?����_����c��&<���S��D K$% 0#"���뚌/]n[k7u#pl4�fQ��#D��s�s�c�fֵ�x(�q1P�HE%HT�eT�@�VYT $@��L|���#ھ��
#� �@�J>3�h���� )	
�"¤�J�lH�)(BD�b��!M%P4`��J���`FD�XVP�Z�q}t>}�{�N����=B-QF���C��Ip醅C}����6ȯRR$;H� YQ11U�A D�C2����������m��0��L>�?G�T��C��������/�����b�=}���g����2QT�?�_tȃ�)����Qj�� �@�r����
 "���Q6�)�@?Av�I��m����k0�⢀�� ����l�Ff�26D�*(��@H&�g����5��faAEAIW�� UA\�2A� �TU9��8�h�F�Ϛ��"_�����d6.����~�����������r��`�j�@cp���ֻ ��M@��TW���*ᤴ��[%�� �74?��<DU���Kת
���m���=�����wTPWpd�6�$` �HQ%$BP�I�$FKs��0�m
@�	���m���[��M)��pE\��"���m��EI@���|�l�.���kY�eU���~|����b"�DMH"�@MB. �U���Ѵ>I@G$D������`}��P�I���¢�$£�������P�B��)�=�����S�g�^j����!�߂�+����E$TAt
?>|��v
���EG v�=8S�*J{��F������	�=ښ1ߙ��RZ��A�#���$M�sw��o�AQ�b��RH[�Io؟3l�����B������	���&��@U�⿮
9���{�T�j"�
<�?���H�4�;��h��/Q��G��>wx^s�@'bA�j�m�{k�c.(}��Ѐ�
�d2�01`��L*b,22@�2Ģ�LB��I00�`�{|�2�l�����T��U��Os*>��� �(rGנ�=0��
�$�T}M�Q�,ʃ���>T;x 'b�3G�����jp���ؠ<�Gt�������������������UG�tv^ʱȲ�0ʣ���A.����C��($�|=T�E��z@��`��G�/`����i�;@p |����m�Oy��aӺ�j��+���Ҩ���=��p���; �i�
C8����
�
;�+�^��U] $�>{l>^
{�S�(����|�|/z�0�QO�O*�G�T臍�@: �>�b�<���4���POTd]��pTwP�b�v�9(�� �ހ�x68�B��
$/�.�0:F ���}.�A_C�����U!{}p
*���.�$ 'hv�����
>0���E8!�p?�x;R=���|�	���xv2�����x�����(&���8<jv��ﺊ �I�'�0@��A.b������=���{L��_�t"+�/���^�XD ���������� �����f{�`����_7�$���T�}��?Wɇ�k�}��_��O���?���y���������/�~�x�C��?��g�������O����o���1)����4#����K_�������E��O7����E�Nc������I�DΘ��W��?��:��o�t�7�O�6o��k���m��*h������?���Ʃ����:�>�@W�ٟ�� �Q������B����X���>�_~@�6v`�6}�	T ���zǯ������C���پ���*���0�	*������
�����o����� ? ���u$T��1 �������M{pС�$�J }O��� �����'CL@$RU�����;*��ޖ�u�p@�?���i@^q�ۛ���@��H(Ȱ�*� �_����vڸ u�<�g�?�^�q�⊡���Ն?�����y1s����S���A��eE�t���p.�� #
!*B�� 2��Ȅ�����>o��~����=;�<��Àpv�������I�׬��Yq;�9�Ύv���c����U�  �>�N?!����+������� 9��*�2����B�#*J�� � ����x��9?�zb����K�?�wJ��M� �svH?���7�~m���w����~�����m������	��W�OX���oѽ5r�U�
#��"Gb� ��0B�����{�����R��'�u���udA�0�b��{ī9���	��~W��gt�U��.��/�>�O�{�,?Ih�$S�J��ƞkOS��VO�Vs`�K���Y4�Q�x��T�B(=�߳����ڧ��C���'�X�9_��%��]"ȓ�����^�QU����)rH�>�?(<�k�WF���zH�
�Xd� ��W0r�B�'���3J��X=��Z����^�L���f������9�#?@�ɂs�3DCF�ϲ�I�0��}��(f֓sv/���{��n1"��?�:QD*@�J�������
U��_�+˭r��� D�=[�
���x�c��_(#� �0�	8�0(m4��d��F"�ɦ��PAe���pҧO%	��;���p��Q�,��Ք!yE��	H�1ߚM����֞�s��S�����' #�1��z���00}�6���@��Z��>#PmZ�T��U�����n�s���'�ƿ��P�-�N��s��y�׮㷫��o��O/���DP�I�I e�dBA�Y$ID�T�	E�HE�8 �_�Hze��h�|B1��B2��'�y��i��&��Zu�+5�`��H�d��
,`>e�=)(=Y�ex(�]y��c_�\Fʒ�Z���_)>P&��YF�Ʌ3u[[4E���&��ZEB�6G�W�|��F����&+�k�M�Ҳ�U<t/@h��Y$���F������+�ޝ#,�"&#�M�M�~,���D��t��V�V�>�x���'�2�Pb쭈>"R���ݫi�����!:���~i�BVvm��%[,��)J�gy�X�V�c�$kiʘ��x��%ZVAV����?O������	,*&^$h��!�q/�ZR��/�����$�hE�Y���Y�O�@85�}�%x��,��ٞ���]��VO���w�j����(g�Z/��;�d\@�վcDv���y�7�bZ������N7V��w]��ZQ���*�v�{M�E��)�+l��ZVĳ�*�mj_�� ��)���z�L�c��z�Z3��q"����)��Dz��E�O��}Z��=�>�\��7��[K��~�]u������ӣ����J�����2� ���=�^��;��紖Z$�"�����AF��Z����4�|mlAYjݩG�K\M�6�Q#�LFoҗ�(�%4��x��i��'�6��&���m�XVq6Y�斅��Q�m/#q��Xg]g�I4��/���]�}�Y�h��M�6̷���ⴂ�Ѷ���c\ѣ���l��v��=�����������a����m���~6�x�� [};*���y�lqqX��7����m�$�/�	D^���Eu�����v|��Eά�s(�[T�M�y�aȳE(����[\�m��i̶#|S2��+��j�39�l����w�Gii�����;��e�8=Ʋ��ݯ��mnw�ѫX���g���c9M�c��i�1D����t��λ�j�����<�Y�)*!�2��z��h��$,z������r7���*|����^]WZx���g$V�z��5N6
5�N��0�
��0�ʌ���$<�'���	�k��f[On�����W̤t������p�>w�δ��[ҭ�ߞ!��\>�㍖��J)�us�j�ٖ���s���Kv۷T�����W�{1$q�:�HqNd5�s�X�i~b!=30�#���0���y�m�]qT�k*	$#}3(Ui�[����_�B��v۝3IQ}�����ųK���ޝv���G�,s��'oZ�g�����=��~�-���� ��*��4"������?_�]��9>r���&I ����{#M�cSWu�[v�Rɖ��́ �f�(�@�D�c3'n<���>���1`�Ʋ�*Y!�Ea7c)X)����
�8�fw
�`0��rjc�� �ǋM9o*c+M�R��tǒ���H-����Ù���� xZ)�R�*���B�4WP�yǪk���w��Zsڞ6鏬�y��[zhr��hᡠ���7�}%����e�H_߾�㦾��an9�6�}��.(������;m�t�q�צ��7m!��>:$�6��(���P�3�=;G�/]{�`����QH��oXv���8���W���z�
Ώ�b�/b���5ۜJυ�y����n�萜u��y���1��nբ�t��:.�۞֣�.�'�{��=F�����c�x;ͯr��m���k���g�b���5��0=ztNQ��Þ��̬ɿ�OIG��J��n7N4^%��B��QI�N�@�~l�M=�8�!E/q���	B���S��+P�T+F<כJ0�u{w�&:��-����t�gZ/fm�'J?]miˮO�s�sȔy2��	���WA����թN�0�@F#�6�ϘŻj����Jڐݸ��>��WK6x㎴�;Z٦q(���_m}�tm')WZ:�)�C9C�-��rv���׼;h�S����9�=��8�o��ץ�f��ě������m��ꃿ^3�:�D���u���w�}�-��u�W��z���<�<�^\XA��3bp�֜�<���W�P<y�+i��&��u|�������t��=|����v��mN���{��30Ќ`��v:��Iff0�m��C+`EM(�!(��
0� � ʒ*��2�@� � 8��f��6͆���>5�=/�Ϸ�%�~?#��Yc��M'^:e��鑾>���Jy߳F�C�v��k��o�v��j�����S��q�=DeM�zc���Z-xτ��nt�n��ɚi��m��{ZZ����X�۪x-�E#KL����^m
�W�ī���9��w٭�Nt�7�������D�g�q�w���^�o�]�篼�m�ϟ����K���}�!�y�ߍa-�x�q���d���J�[���Fv��-!��o>���1��N�4�ھ��׎{{2�O#�������2��}��9j�����Ӈ��e���=;v��[sף�m9�X�<��?S�m��޻��MT�^7�o�۱n��m*W-��Pw5U�}s� wtV���yqmBJAH���z�x�>�5��/��N��_�ž>9���������_׺C�+�i}������bQ�v��>+��g���4���m���O��n4����u���7�x�Q��];v��8�~�Ε޻w��v�ޣ�g�`��u�I�4�ײB}���5d׋��o�����/s�����t�������Ϗ�4�e۬.q�=}�o!���p�ҝ<����q��'O}�'n�%�=��w��hOsũ$�qC��:Y���xm=��{��:��>���^���O�״��H5��v��i?n��ic���e�뼄��_/��S��/�����ae���0�����%�_I�҂�k?o~���N��~�[�Ƽ&ͷ�'��l�~��G�>�ś�� 9�}{�RQ��T�?��=W]��Ϗ����o��Dǜ���.��w��|���cړl?�ǿ��Ǫ����E�U%�v��h�����k��w����iN�^|��_�y;oc��q�]��yk|O^o�4�=��~q�i�;{{c�	�O��>6���}�X�
������ǟX�s,kھ�?��Fu�?��#O~���>:{�V���!�t�K&���zo�gW��Kߎۿ�e����m��m5�ǲ}/�񜝆ђ�����>�x�-�j�˞~={'���E��PI*(�q�(�]����Xr�-!Y}GYm�!qإh�Ci[�w������p���W������c��+��3jmVPԞ3� �Sc2�X�0S�,��D���e%���%���KQ%B��"�6�y�	�	İ��sRr���n@��$�d8y�83�P�"vP>)�NU@:D����ӷ����4��Io��֔�߷������>�:��<���okkߡ۞��Z��N��������Ͻ�t�����߇��8>����~o����~'���Rx���|*�_yw嬄��Ǐ����B��^ܿ|S�u�j��Oy�㿋��2Y��~�������hm)6�����3�o@�ިԺn:�}���*[��z�G��O��_=�|��u���5׿�����h=Z-NG���m}v��v��~����;W�~b(Ю3�u�zm���8���o}�,<��~e#�;�,)��ӏY�|}`6�4��6e�c,/��8� l�:Qp�B�B#$�m�t*�4P��K�~�Yt_a�#�t����-~z��wޞ���%���+hs��|}���>\���/o�W���>���q��m1�����exD�^6u�P��"W-���vGMKy�f���rdBq�����b?���{Pʽ���}m�3��Ӫ#�-�f�|�[���������]��0�T9u_�
h�]Ǝu�D�'|�X��]uHF|��х�)��ao��:a|i�	Px����y��&����� �	�GIޓ��1x�{f<J����*��AQ���@��\㢼,�Q3m�Ӑ1��X�#���̱M��n��Q5�S��a����r��}�ٔO��_��p� ���\�g!Q�iR"�C�E*�?-6��>�mDt0���� �$C�����s�7$b�e\�YvP�؜�IC�2*KL��:I�!�%�(E��.�!���Rm�Y-�h
��#�	 �
c*F�L�(��
nBl�2A��d�2*���ʂ���K1��L�e@sǺ�K$�Ӆ8�e��uX��'f7D��V�D�dS䌴�d�d�X�4�D�J�!X�Q�����v���������^5�b�o�/]~��v��A1�1�4	�
�9��Z��tE�ErJ�Ûf�=�G]}���,�)ӈkJ����Y��vS��h����s����H�!�Q��!	�Ŕ�D����.F���Z����Ncr)�=9�Z[����8����ό�n���鼆���;��Ґѻz_��ȟq�;~-ڍ����O�*��ټO�W7��J������)�lP��(�SS���#��hJ�=<QЛ��ydh�p;�Q��a�g,�ٜ��\�F�c�:��JJ9��%@�^}H�xG"/ 16ǁqRM����+�>��v�4?�~��_�Y�Uѿ1��S���a����Q>��6��Y�/�c�Ã��O��>:�b������Z�TzZh9By� .j�ȕ<JZ4����HZ�*�梈��Q��&��Ae"�H6K���� q�9�X�S-�0������c��+��!8�U5YI���_1�U�b^�TG"e%>u-�"�[��n�*�D��:�I�������p�P������G	3�Ȩɐ"�jO�kD�o=!e�ɂ�R��V*2[,'(��s���Q�l�͌UT�B�RZX����jR�"�p
��H��
�ʁ�i��8�EI(�(��p�$��`��J��@�2(�9(%4l�Q���ZD)��;)��`Xh�.d�9`���31��%�P���5VvUH���LG&f�*� �R,�P@�j�7ȭ�cVqfi��zÚm5"b1%}�X0L���͠(6Z
�QɄ	@d�MY���EY���1o	�U8��L2�\�%K��H�h��dUKBG��E$ �La�(\J�\nMe��!�FTwbv�e] ���Rea˙y�=�̀��u��5�^��ǅf��U>!��
���=�Ju��B��n&� ��K*���c��A�4�b��("���UA�<�E��LA$L��-�\I@��f�b�i'�ؗ]&Umh$Ӝ�T�&��!��I�Jx��U��	8�̔*6X���G�L�Hqᢟ
@a�u��	�I0�0UȤ�����w��I��qĂ: �u[J��M�-�D)���e��� ��p�ȘS ��j�y��m��͚hDhJ��+x��E�� �ӡ�Z$�8�Rx�M�^*E�����F�l @�QC�X�"�["�SOKV�Wh��P��fe[\de-"�a��`	6�X+���Y��)�b.��n3kȲ�5X��4��q�MA��y�>��Z� �����E�^iG�����t���1��H�[�(Ul��D+#R$A,(�(��R��~THnD��Y��4��v�FѱSP�h����c��gG���=�������?������}~�p� ���s�\����@��@�� B$�2,��)*J� �\� x���|����g��~��K��}��=~��1�'%���g�Uq�Z��aʨ�ލ�O�˫���ڛ��
�9
��aE)U`&U��i� ��Z���D�..��9�Cc�MH a{����&\1ʅ�Bu���Oy��ͯ��v�x��;�F;��6��5Q <��Zd-X+�� @.�;�=bII��Kbj�*Tc�~�AZ�URҞ�����Q�D��9�@�����zg��"��Ʃ��c���@7\,��V�b��(d�	�* B���a"-c�l�'çibi������4�.٢ -B�|����/!d�M����˃�Ivb}Òt��
i���$0E�~����ePdRM7
�8�j&'��gYAB�+hV2�r�2����O*��5`dwk�FT-CF�n�.f*�*SX���@�Kb��T�E;l^�����n��a�I�1Q2<���O*%U˗���4�_Qd�%G�E]�*�vJ���I��\�����T��A56��"�.��,Ek���nA@�+E�pc��n9�V�0��i96�Z�n�gA���u�,�E)�Z�����J&t��)E��H�>*��k�Q
��&�.F�9��W��� �X8�L�R�0�����44�x&J�z�l:,F�8�1�
d��U��0��J��$$L��h�8��TW#|ԬR�׉h�p �������Q��*�l�*�1�"L���Qcm��1VY$��`u�ؙ
�f��l���tu��T��ԫ��]�?@#��)2�N��X�*z��i�yHMJVL�lF[e��D�Qs;l����=0EщL��X���0nj�d�g��Z�H�F����s��JIEY��R�=�[qW��6\���# �Ldk4Hʹ7R��F �j�r��� �8TpQ
T���F�S�D �L��	L6��5��y��YM_O�%Z�4�"�"y�
��IA��*�Bj��FW��P�J]peƀ��9�E�ځ�X(�-":�'�@��k�yX��Y�V��6Ԙp�G�=����Y�Þ2��J���TI���NAK�RQ�3�1I�M+1C8��}}}}}6���d:��&CG�����K�e��[g")��'r3eH�k5�E-�V!��&�|������r��Қ�ICs᐀�6ZJ�PO�9���O,�c�Z.e�O�&���v�o���?����G�����t��v��o�c8�}U!\^�Ǐ��0~g
��d}UR��M71���Z��z�1���!}�-�m/�8�j(�Цd܂L,��]Zx�
a:͂Uc:a�eF�b���u�
Am7C�9h^JWCU��D{�+'�)#4W<g�a�*�J^�.M�P�֛�`F��G�X�ѡR��$J�)�N�"@�2���䨄�`Hz�����Ι��B��&�նAe�1�$�0,sL0�)��mD�a��B�aӳ\���Q�j�`����m����8��э$����U P����C�,R.ف�>���#�R���bR��s�%��5b���ZJ�}!8�Ƒ������ '!rDDS���yI���:%N����
�`&[Zvs�-���(�Rٓ�d�iۜr�k:������&W������u��iX���5�$+T��P�1T��=��z������f�$A��UɦYq�&
��d��|"�6N�Cc#�]���.��p��ű��NI�@���n�ǅ[G�w�H����M5����U#
�<UGz�7��NY��U@�A�Z�0bR�8%�Tצ^$X��N��Ԑv�"�GX��"  �`�@�2d��`��*R�8���)�\�h`�%��స� ҝ� ��H�&�9@��#�$ �
�C��� jjӎ+6}C5��^���0�@�0�$�Q�8kKJ��k:�Qs:Obfo ښ}GxQ�QBD��l�T��]�����
�o�Mq��i.�l�hJ�b�Z<Ԝ<w�1�Zl�;�^�hQ�>�#�A�)��0MW&�1�D��UhJ��fl�C��J8�(��S*T�$�lٙ]�ˡ2�q�3FR����6�_��<|Hu�L�єIF�˒�+l����D�6����J&���@O�M�Y:r����(
˯5)c�����0�sE�Wť�M�Mmx�B��LH�S�B��,}��?�8�L���z�+ �f:+����Y���v�T)���#�P6mf�CO���I<��,H��f��1��Z
�4�늴m�g�\�H-q�Ƅѡ'�x�
q��,Y�
�#�̠ � }}lŸ�Hn�i���E��=�����n���S�
Q�(m��;fƉKu�$7-!W"�u-�2Z\���_��fk/�uIbf��PMi���nf�-�dѝƔBӊa�6�G	K�),DBx��!ш]�sew�z���*%����ԁ#cj̮�#A����k:�#So�5��#ʡŕ�M3jM�L )�T_8��"�K8�N ��u�el4@�aK^2�1(�e��x\���˓�Y�x�i�7�8�>ZADf��d��4�D����V�܍;�_]ݵ�ʴ��Gi�� /"�P�f����w�{<�����Q���{�v[�d���w�?7Y�ũGA��6B)R-�" 䈑��ʚnm��l���.
1�.e
IFk��F��9�q�U�(]jd��cK�cr�4úLQP�	�"HOfv����nS�9M��ȉ����E8Q�Ek0mv��E,�����W\�|�Y�^5ڝ��=5[ZF[d�w)�t��w!j�"x�7,I�|�)8�I����.��n�Ii�L9��p�M����[��ϞyԈm'cr,����cF���S�v���pgr�+V�!^KG��Wd�FI�)�.zڷ.A���p�J3 �̞�@`:�=�<���3�+�,N�i�~<5��#|!<u(z=�74E�x��^��y�#a�������	�[-�m��LWO j^��V�M��}g���3Yy�X����ۛ`U{B��PP� e��h�xR,�9+Y�(*�����E	&��l��,�E�f�m���1�2Ln:($r�� �aڌ'P�# 3�Ɠ'���y��d�X.��/>���'v�M@lq�#�e���Х%�@�M�U5�W�	�Y� �yp�n4U&
B�y�-ő����9�z��&3'|'ʴ4�<D�����0xp~k$x��]c=
�Ht�e{�]��~Q�YG��%�{K�1oai����[G�v���zt�!h�kG�<�f<��K��YN��CsՊZ=jv1D����}ciLu���* 7�j&��3OMt	���ε�M��a^���hP�	qePZQyD1y^a�O_f�����	Ee1����TĹ�9��YoE�9�
�;�o62�}�4%�˜Ҭ�m�1�#���ژl�fev�>�MԚ��"�i��[;EUaVD0|e.Z�R`7z�rNr>�z��Y�qK��1��5���q�B�sx��+B2�:B+��2j%��<D����,C*�_��r�2@�twRSU�VO�}(�0�B��=��Y����U]
��F����@ h(W&�"���5�Z�ҵV���]o6��Cԓ���Z�$&� P&M��Ia,\�B0+,�`R'�bE[R���@L2�s,+Q��[��:��y}`���Ff<��K��Z@�_����üJ J�$��(�J�D�@ �Q
�DA(Q(D�Ph V��PhR� �D�ZDV�DJUJ
TD
�JR�@�EhD(@T�Q�?A1��ѵ��3�-�0�V[0@��u�]�7 SDo�Ӗ�ؑ��(hT)�
)D�ɠ���!>8	��`N����/v��#����������=ϭ?��#�� y�D��J%��%MI���$Z&e_ϒ�E2�,�H�E,����@�c����"D0�S�]��o}��b��`lBP�R!�T�Xk r(G!Ԏ�v��MJ� j!�v�$�1
[0,�
�$rWP/����xH�7�8B��DԪd�$^_G���Kϑ̳y�w�|˼��]��y/���n����@8�4���h�5 ��"c�6$w����P��MB<!xB#,�
M� ud!� �� �wwШ�d��+}�5(p�v�R�p�|�����
䦪��[F"�"�@H)��F������@;B���*P	�@u��yL�B)�
�@74b���&q�x0�Y% �7�Y〦�R�H
p�w 8B�� `fYU`�,�:��4�(���*c���悱T�0�� � S3xW%Ӊ��٤T ��M�2Eu(D d&�(� 5ƋF�ZE9B�v6-hZx@+�i�6�%h �P� ��H�B�
d�@��±PԢ�,E��@m$JZ� �L�N�b#�h6�B�J�rMB� o*�J ha0�MB�.�rC`H?���H�}O�{�O輷��?�����D~o���c��㾿4��S�drT�c�_�l���$i���ˊ"%����.�D�~�㉄�m��/�XemKQ-�l/Ƣ���?�8�%%�w�;� N}d�m!h\)���
��1�0VL�:�������`��l�f�Uk�a�h�\.c�j���D#�H����0T��`��h7lt��YE�/���Iơ�'y
�R�A�<�c���ji!�Y���3_'�[XAx.T{�β�Ջ�j���I �|
�DR$E6QRNMe{B�be�k�$�
����}��_ܳ{�N☛}�ol� ���XN��<�i.N�届`��H�Lǈ�(��)53����7���y�v[�(�e�S��У! eU*B��P�Dp��o��IQ
�(��o���	Y1&�]qh�^I����k����&��箿4�|�E�w*~,�_e0���Ǧ��3H=C�ƴ	�,�w(�Rޞ�e�@p�����.���{�5�r��NX�>a�g6:�v����f�V�(�d�/SNԷ��1J#"���P���䭥���di�F0{e�F*��#E� �e���C�Y�ӧ,1��Iv���m��e0�4�c���*P��&j���-��~�L��]m��4٦� Ҏt� �����Rn�u8y�m��`��؉�t� �r�۳�m~���E�m$$v����,��%�/+�\�TԲL��"���P:�m��-��P���x��A�3���'�a��6��Y5�I�$M�Wvp?$�\�f�ړ�����l^Y�Ku��ig�:uS�~|	���`��U���-x�ԩo��ފgKa6r5.&�4	�M&S�����}����e�� �&�$a5����Y���v�#	:j��`:+C-��� ��Hʐ^"�@�B�ܛI�W!d�.	1�M�(�*U*|�)�����P��KIb��P�9s��N���z�@�L<�<1볃�_6��k���j��0�`�������rS�������!]%o0��dv)�{4��u��riD��L�8�^�Tr ��f�����8�
&)��e�M�"��ydA� �G��!MŹDD�Sm7fD��9Q#��}�����ǈ7v{H9)H��R�"��-�=��w�\��D��<�x]�{��ƜĂ�9�.@9��ķ���!�I`�]��8ǂr�qk'�;�j36�I�wDqBn*5�OT������%*�bP@����`��p)���e�s)H�j;��J>�ET���Ne(�B&�D�!�Dm҃ ���Q����7bUM�&	�@uZW�a��'3���9CQ$�b��J&��S#<�X��)p�41 �l�Bڌ&�͔�Wx�m18!����?�k�թӬ���|�>��;�Unr���E�f��v�I4@����`�_�@��F$�~��>�~��7��>��-)��TP%V�A�B*��P(�P
P�@�J�9" &@*
��T(P�r��D5�� ��W�QV� 2]��D�aCh �Ti J>rT�QT�v��{��oC=wXTiH9�>����L�)�\?d��G��D~%g�X�B'�J
�	jA�KM0��Y:���j�2�P�B7���h�J%B�@̺�k̫�i:FJ�)��:e�4Yac%�D��Vk��>yH�<�.s9Hš�5�J��\�V�x9�)�$����F�G�WY����=�R�X,elA�h�dRX�[�4���ű��^����5�EVz��DadW���d�Z��4�dU�p�bVM�Nu�B�R�1�a8Y锼�9�)��ލ!v�D�Z^�B!Q9���%�e<0ҿ�*�H|p��|h���d�Md �T�y�������������������������������������=(8U�P�@��^3  �                                             	�              P=�               J �B#L�B��L1�     3���,   �H����($rQ��TIRR�)"D�DH�$D"	A%�x         �z��         @0     @  !        �x  p      9*�P�p    g      �@:�     \ p                                                            ���     � 9�      ���O��E�    (                                    �                        s�  |z ���ZS�m=(@��  H 	     }  ف�IK    ̀�� ���P   @         ��"    8   �}0UO       �I ��4��b��O@h��=OA�d�L�44Ѧ���� 4Ѡѣ�i�2i��j<�CL�1�Pjz @��Q6M'�x���4z����b�����L�z�=!�� � �a ɑ�`0�0�S��ХT��hz��@��    �    # �   �&     ��  y�J�L��5�L	�FL&#`L  0��a20` L0  �� �	�  ��)$ ��L�Hh@ ���     �          �    ��@B �dM4S򙦦4�M&2a��4LГɣ)���z���5O�?G�S�O�O�=2��jl��'�y��5=OSM=7�jf�$x�	�����\�`q�5�)�LdTX���֗k,�#��~~�\�������	71����N���vu�VىfVpƌ5�
#���Ԩ��S�^�^�?����u���&sIq�c���ڶ5V��f�Z�[Y*��""��۟wTDTȰ�֜����?9�J��&���w�}�Fj�"�T�,�5�_���x��}��pE:�� ������:yI�V���VD��o�u��[ �!�0D<�?���m:������cu�V�f�j�n�v������k�E �24��I�:N�����a��+fTV��
�DBI �?{`8W��U��ȋ� ����̥�5s��C��7�Df�4�ad�#�3-2?2	 ���8� �&�Dt뼁cU����E[����h�.��뤆 �6z˱�u����]w~��%5�'���x�n��@d7+j�5��[����L۵���s����u�`ו��L�ѳ�1r�C���bB���~�鱌 B��3��~�!5@�t�h�WM0������b���a�!�P��=Y���W�!0--�,\��2ʰ&j��L�V�U�)e9�"b��"�#�$��sڇ}��#c�������\�Ukųxy[��׉���S��VchF����p��a9��+�=0_�|�B��)�j�𺆄�%%u`��0Ĝ�ڬ�$�AeG�l��S��cAZ2����E�N|�1�ceVr�Q�8Z"���KXzK}^�)��̈́v�[���C$f�����Mm۸����"#�����ӦZ�]@"@�܅0��p��\�ll,�Fd�ڸ9�˘���-�:����Y��К'�[���!	In�&�s�v!$h8��p7D��.��U�ゝ�NB3��[v>Sݏj�>�g��$�����?=�af�����z�@l2��ǫ�EE|OH~���]���;�H���Id
�%�@%�1�FF!WVk��5v�J]�6I��$����pB%�r)��3�mV�욖l�d��"���E��N�/A�	�+�� �/X�*��&%���wnb��m��.�ru݈DВ�n����+��Pӻ�Hݐ��:Q9wv�w#MITD�N�A<�E_��T�H| Bq�b��F�IX�i�b4���B)w�*�����E:�$(J�(*���)ʌ� �),�J(L�R(�F����;ὡ?�ǛnG���\��0�u�P�$�B� B�	 �H�$ �"��¤ D�G���7(��-� ���{������a��c$���{ۿ�s��w."���ʼ�[�{����>?��]������_%�������{c�^7�z�c�������k�~���׻�?������y�!�ގ�}���3�z�|Z����e�a�e�lV�P�m���O�~��*_����~��|���w�Ay��~M���~�?h���F ���ZD�	P|�A�����qO)FO�>�>=`d	�Fa����}$��C$@=��66�^���q������l߇�G~<w�>��N�7����|��<#�N�O�v;]�x@T9�L89Ç89���zN��K[���/����8%ҝ'�u���O����<;� ~~맡<>s��Ps����DTP�QT E_����������i�pps��?{x����{�U�	�����w#�+^��f�j�G[v�z�R�/�"@;]S���d�D�������֫-�7Z��)(����k����N���a��9��Y"� �vF��h~^��d>���� ����~V>놠�b"v��U��l9��߽�9���ZugG���w|��N�AS�~|�m�sp�:��տ��*#��8w��6ծ[* گU���{~�o��}c�G  �{�[�3�=�ٹ_��i3�Yps��>P΢��*g�^|W�W8:a���?�����>4s���o�흅)��s����)�� 89�w�=���ו� �������<�� s��Qx�]�9H?o�����l; �ps����{�g���8;��ھ�P�W�9�.s���t����)ky� 9�9z확�"�����?t0 γ��N���(f� �M��K�������?}|~�{88 �i3տ}FA�ps���9�nV����P9��������, <�㉇ ά}�u꩚<�N��s��}(��G�G����}]=�C3�����pt �q�mի�U�xw��O�nwU���}K�?�9� 9�������>vթ�#�A��t�m�9������޿w����� ps�˳[��>�����s�KR�KÍC�� oߨm��!���~������3�� pv[�'����� p��z|VGԟ�`9ݕ�v�r���͎����pp��u4�.a��8;�'���?ZJU�=� s�����P��ec:�Yg���e\ ��@�7�n��P��MJ��� ��6�y���8Ag�ږ[o�����[]����>���=N`89����Ƚ�'��o��������uxp�޷��^�yX����pp�G�I�&��vn�s� s��\��I�vwŀpps�V�<89�;ʿ)X_�
  �ox�*����;llz}k^�$
��w�������z�lm�� ��hĭ���ZV� �8���T��AT��q+���6�YD^��8�P�V�M�*!Ƅc��H�.:�B@��L%A��K
0�;�֬d+r��U|4�i��C��`hE���U�|OJF�@���+����	�����I+���Sθ
6ާ6˖ @�	=���G������O3��V|�n�5��kZ��'�RZ�s���z Ms�rbB�}8��|Ə�qM^i����K��I���ؚ�c��H�}e;шh�}��1H��,	@��`v�ܧq<ZA4�z��]�z�zV�.�i!D��{ώ x���z��5���v����2���u�Ա��/l7JB^��Ҧ�](�|��:e�k����HV@������U������fi�J���H��*���y�	�LH�x�qcY�[Em�����"�<U��!R�˼���,%u��Z��N�]`@!r�@�fօpT���W� Sͧ�B�d��20����r>��G��m���K-K�m32yy�'�I.-�mVW�`��-;v�ZG�j��Q���ǎ�����s[j��s�,�ԅ�k)(�)��@�<���ѡK��@.���e/9Y V���qb�^=
\R�ำ>,��9�/�EQ���"t"v�̠�x������U�VU�̞̰�yJw����� H%���ׁyH�YG�%8 kd9��'	��yHy��r�Hy��<�Ra��۳���/���)<޾���ޚ��6Um%T��>{���[u���[S��%S���&Fb�(3=I�ȉ�3�(^ᔤ����jj���+C�<���-b$�x@��:c�s��z0#7�x��M��ok�%�< f3ޗ���̀f{%(�&��2���'���
��$ş<�m���@Η�I�"_6{K<$Ozx�$x�,��*�'�m�"���g�`�|_̵���= 
��aX L^��moxQ&�O1��POFᘄ)��bF��-�c��f��z�t	Є���[��_`���M�y
ߺ鸐u�k�N�����oJŶ]ZAI]RM_]*F"AP����RQơ�yf=l-��Q2q�Z�E�v���BA��6VG������+�Ӓ@��ob_:6P������Yb�&���]��a3��S�g��ix�;޷E這�	Cl���d�.� X2$g�yTR)�mO_ZP��>�Ϭ�����W�Kր^��Y�i�[O6�ޔҗ����U��8�0F�i[�V��6it����,����K֓�ͩ))	R1<7b��};������.X�H�}d��'j�zy��<scB�85I�P��g�����3�/��:�8 �x�Xմp��P��m�cĞ8���112�-3)d��_y��:�{{r�B���Y�Z�Z$�\nRz�)�UW�Gy�!������xy@���z�6Cy�e�b�ROb�����Oy�OF�M��B�PQ��W�Y����L0��, ��|_k2Ş��|Jk��'+�】�,`"�<��3�
f�����1�}���v1N4�Z=������_k����vP�asA�4UUBH�B��v���+��q��_:�l2�{R�x� (��}mS���$���п^�!b�@Wũs�C�k6~-������J���
0��k ���!$ՠtkc�3n����@
�c���x�����N�Ĳ��N��� O)JD!�T<u���Z����Q��l���eű&��a��@�D�'�t�a.�x	��ۼxK_��3@�S�L���������4��̔�ӾO�Y�~1c�
Ie勎�a�yc	�֢R�@�,SJNu�&����֭���>q���j��o�$�I�� �"�zo[H���l�)"R��}��l}	)���%)�@��ʶ�ڐ2�|N�t+�z]|q9jD��z�����B�֒��T	JR��"	#�$HKm��4HG\R9<ڑ"��a��Y�%��i�� x�z��|Fd��I�4���Ǒ�!W�BZ�QԀV'�Ӕ�ľ��_wt��F��<_Ho�����B��ӷ[��[n���ߑ��wH����aW�BܥckX&�t�%�K�x	VY�~�p� ��*�Zڢ���tĭ�!!	<1d����!X!T*,h#"z��2�,�m:�z�ŏ������Ğ0��A��L�,�� 6ƴ����x��{ 9�I�z�Cվ$�P��}t��{w��V����(��l�a�z�d(Z�yp��ule�<zy���\�J1�)�Y�0�$u��|	�&'C�!H:��� Z;kk�����'��4��:cSlX>��Ď�}}Ԙy!�`0[)2�m��A��,OĘ�`P@��[,�/Ke"�)�2��E�JD7mJj�Y� ���q�ֵ�C���'xNI���bb� J@"�b�� �:���K�%F1,%�-��,�X1�( �\G�|u-|Y�ՃD�-�g�I�z�{K�S���B���u�/:]���Z+Z^%�"NNlYb�/y�X5����KUn�$���� J���ҳiOb�kf-d@N��KU@� J1S	Ǟ���O24�߄������4\�H����Ri�Q$����#u��Z�Ћ�"D0�pR9��x�N DzA�l(�9\X/���qh��|�y���|��fO����z)�D�J��W�y����'�jO�N���H8N�6�v0��y`�"�LA`H%�D��Ы�H��(�֐��k���YM,�$�C�`}����7�m!*�'̚�HUU�Ç�+H��lkH�@H���t���� \�$�Ƙ zz<G0�YRp�9E`S��g���U	o4�Ĭ�R4Bk#�Ņ��e�!
F6�QAg��V��K]�	�(f�T��Y
�|0!U;�C��z޶R�U�(��km�'�7�hu� �jK~��ҒC��	!$	�N������8��e �y��N��|	k��KmX�X������K4{�䫐5��:�i�)D��6ZF���X�O/e�M�i[��Y,
�l� ޺`�� 9o0V$��Е��GA�֓-f��r���A	��a��Sq-\���=bOQ�'�\Z�ל�yH�O�I�\i��>z>��WŒ�=[ޭOA� �HZ���17�	�r@��D1��ާ��0!!/$b��-��a!em&9��P���f� ��kIKZٛc+?R�LD�||{8�xN��|HAɐ��aW-����L��t>uBy�-MiD��)
�p+����� ��u�g������\4r�>ii�:�MP	H� �xy�{YK�l�s6������7�����e������6�k�ϟ< K��K���[H4���ħR�V��!�15��a�����O �x�<&[�n��$�:[	Z�d�0O/�(T<�_24f)eH�ļ��a�$@������KI�W�<!/��!�m'�J�-X���3%�N�����+���P�q���,�`�P���cҰ"ul���@��F��>-IIHC5�NK��$8�%����Od4I����gЍQR�OYޯzzy�$	�ybmq�s{\I��혓�z_0��@�D8YYnn�W����9"0��io+ȱH<,��N�-�__1za&ae
��KYeQ��E����@<�u�D��(�^�H����0W��Xg6P<3j�"bk�f�"H(�-�)ذ�}R�	E�q�&9)űDi�8 F�q�b��1I�0X��x����2׽��O:�|z�K��I�Ŷ��H�����(����=�͕$@�
JX%o�5Bf�h���
�Z��b��P��a�g�J�ĥ�+!�ٳ3�����Ў��3�$�����-��hG�!>�
H�>�ix�RR�x�}g�ŌJ�x�RR$Ƽ�Z��b&#�&���%PЀ�0ԐLZ�C����`D	�!-eRy��%R ����Z���Ę����<��hA��[�6"Ey"H�j�(FVD E�$Eg���=^� ,q/HE�4��"O-C�S����,���@��@��)(���rc��H�^��F�0U�X��JO,<����D�}y�)¢$���k7�`	�����LIe���<������3ꐅyb[#�D���g�0����V0 !��̥TG��a�JMY�6�|�'�Ia"N!�:����{Ƅ�%���D!����� 0Wz>8)�{6LS�X)������h�-! ���uQH�`0}R����x�����i4@��i,!f�=�&�͑$k$2�-�x'0C�R @����ĳ���,�R���f������r�����.�L��X��О=+0�K���B� ���"q0�Y�	���=i6"����ے!(��c�:	QQ[B�*���R�1"q<�#Q)�(��*ǡ�d��yV��a�&����(Z�Q,�ByB�HxŁ���ie��!���XO2�I<�'x�[�;�� q/��׆R�o�b�9$s����N�aIf�Զ�K������'�T�0�_�� �g������`VԄh��1,������!1XU�z3̈́�*�.3��/Ym�0#Ƿj��o{`%��z���0��J��@�#4�����=��$3�.���e�x��R�e1!lHXV !�-� �9|3/yp����y� #�#X�H�CD
�����ա+%'�<!ʾC���:ڲ�ڄk�:�	Q���R6��Nb���R����z�̅�uk	��m�2e!�Z�d��hu!��x���H��,�[�_VZ�&n��J�"����� @U������#�UszR%X�Ky�V8��UD�S��m����3��i[-��"q�vR�ϋ�!'�/���16[��R�(@�Z�Ƽ1P�B�u9��R��5��G���%#OX�[zSGz�h���#e�����2�,�	��6�HŦ;3���[��d���!�!�+����xyZ4�ԩbȃ��.���#%^���z�W��5�@�%��IF|��=3�GmL����捑"YX��T!�+k>/5�M���ן7�y����Ov��<��\�bD#�z���\u�B����!���d:X2+��&�ƶ���!7�Ő!��@m�(��2�٤^'�t`�͛����z� � ��%�OW��"Y��%-��C�����JE��K�!"<O)<��(;i{Bj{P��t�c HL��\yh�:�$�,��F��5btK
�e�U@C�B(��&9�X���@^�FǴѤ'D�3ڤ�*�+-����"bFJ�-e�>�u͢�S�
K��e=Y�@
X�IHm���f{`� ���u���s,Js笇o>�%�q�l�ׂ�޳�B�u�
�2��>JӭIF�HX�(e�`��4�{������2�d��R$��8�^X��(0�Ұ������X��w��O �����Z^��A^�� j��s4B){y6�����4�'�qd%`��5a����{�ޱ�b��I�:{�/o��A���ۦ#cx$%X�-aA��(_>�<�k�@�	�K*CJ��zɈݺ�	3F��8� ""B-a ��J����1�=�z��/���0x�V0`�f�Vס�9�@�j���p���m�{@���g�贒�6�Vz�ᚩNH�,$XĈ���lV��K�1��%���=3�fx@*�{�gb�@�;3Vb��Uy�3د�U�P	�J�D�@�z����A�R��b>:%X����
�z�ۮ�gX�%Yԓī��`�y
L�fj^�	�m�9� �Jb�T������2i z�2��4�i
��QE�j� p���hpq�u}e�}�=+>bK���U����D��f�[�%�:�o-:�{ȶ�J@-���6���H���٘�ty�p��<B�Z�$j���䪬<M�$����Z��C�g�uMAR�������WgǬIx"=GX0_�V1���h�f�����է	%e+[}�s�����s S�Ʊ�<t�e1��>�
�Il�Yf���+=y;���!<M� ���WŦ�� łN,�&̚�\hOi����g���� �V�����i6���1�y1E��DakHD�Wϋ�q�#X�bB0�l�D1�)�	���4A'��Hy�R$ڴ�1L0%��AR��T8�&f�Ĥ�Q��b���l���P!�X)/��Oy�)�<���$�$�����؜�Y���y� H�Q@�		Rq ��[�������������[������5��_��q�����E�������� f������Q"��}���������������F�s��G���u?�U�
�^�H���o���G���'���{�;�{|>������c���� ���&�?.鱮)����:͟�����L��w?�Jo/+o�3�+�PM��o�I�X��opNoK��^��D�j��0��d{H�E�e����W���׈�h����� ǀ|  �a ������ 0   ��g���sü��מo�W3�1�9�v������8�W��?<-�|g�M�C����&k�C.=3��)��kS\����ȥ=:m�gBd�&�F�U�<��4��K!�٤���w�JUS)�L�V����
@������}�h'�D�b�;4���	��9��{��a�s�]�����nv`����K�8ӻ-�!���i~VCn���vn�3��w�ׁT�Sf�S8L��3�E5N�J�V���t��\S�~�-bz!����V���v��Hvl�M� !�L�9#��t8�}�GI,�@�ç4l@궱a���y���
q�Wxu���f�E�/I��cxE��DUD>FE��NSA�lJ��OCv�U�1��D��- �,���=9inW�k'��'5|��C/�m�œIӓI%RK�m>��9�\�JO1�@���0f6�	,'h�X�)�d�ի���jݠ�4�"K.�Dё��.ܯ&Xa��VS9+���;Э���2�}�w�c���������l��G�4�&Ք��]�����ā��85�s�9ew1�K���$g!�;S������i�J�
��rƨ6?[��=���qOI��Vwl4p˨�&�/�ձ���!�c��D����3?�c��1�܏9��N�t���<`��.*S�3R��QW(!A�Y�Q	3�O��r!�� ���4l��g��4��~����D��	����n���@�|�%rN���,�<�d3D��q�� J��'p0-y�χd^z��^KIm+�?=��k��#�����ȪO�yt�v_FC��ڨ4��A(�fg��ȋ��zz���}g���u��H�'��T�Y��!�&n�6�.AH�1��;h�`���;��j�4�$�O�,�F�)�Pe��w��������<�r=U�*X��4xC�\p�^�1C�4m�*��'�F����\}@fCV�z_S̼�ީ�o�O��k�P���Q��;�m�6��;t<��M�%�grJ�i֤Ā�J����3Q.���c��ø��.�n��,�{�Ƨb}�Z���^��SZ�k,(�b�#���'���!��	��W�.3��U�![�Z�����;�Z�hS;2�n�oK�v;�����#5�>����j�N��Ҏf#}�z#�"�|XF�Z�oU�@�v�R�D6��¹p�䬆�ْ��^y��vH��n���x@��r���nlyyȷ�x����ԟ��R�ەBN�����U����4[�Ry��"ܚ�M�S�x�/(�i][� ��b<�������_i���,�Ծ<jB譪���b�Q�&�j�`��N��R��F��!Pb|��҆e�l��ƆAL� �����ƚ���ͅo#��u
��ϲ+[�S�VG.J'���$�M�O!����ޖ�����P1�+����rq��P5�;T���b�b��Rꄈ괱��q�8����"@�I�A	�O�f^DYĜ�.ĸ����   ����%�	P Y�	~� `��E�$/������3������3���~o��)��$���_����� f��o����?��С�1/�{�X9�X��?�	uH��>��F����?��#�o�v���S�EN.W�J�_�9d?����7��ؙG�L��9_�8��W�G���a��Ĝ5����g���e����t�lܧ��^�YLvK��,by5�'�(�W���_����S+��>���"ш�dl�E�(�Y��z�]ڐf����NGף���S?D�RaB#�!�x��BF��;Ҕ�Z��ތ9�����I����[i����9�z��B�@<���fKt�jQ��.=���B�8J2����|���B�m��Ndr��&�1i�~4���6�7To�⌅�6�P��s��{�ߨf_�e�v�_�5RPO&|hGkk��U�+3�rr�#=�X���<��-���'�Y�H����b/i��:�9�iRq�ڀ��2�ɻ�_���P�"ߐǣ6�������ӌDG�^q�~�-��]��[�{h�T/hu�|�̅�,��#���9�@�)\��eV���G*��(l4Xe�h��(t1x�m�}��ae��9w�Z���f(*��B�H9��&��5�-��'�o]Z���a:���V� q-�>�H�2�|K�(,	8����zqy�҅!;�քv�ŖݼNw�u��ҋ�%"Ś�]	����z�>X�֮iH��	�Jɺ�@��r����ߺGxi���<�@�߂o��t��F��\_���lB푲��P,׈�ƞ�>z�;�d˽CL��������=H_V��C�>��4�
2l��:[l���˚�����$�,y)^����T�ĊȔ��y#J^�j$��d���XI�tA+���$=(M"U��J�!H�����.�tPb���(�
�J�Gu�	� ���9d�+�-eD�E�Ɲ㸒W�{+l_Jg�R�]k����58}H�~�$�y��eM(�+)
����>Rn�ţ�u����bWr Y���������r2c��SsE�N�h(t���<�� ���"�a�J�>B}�L0�|"�𚈆I���,N�T/����Cw{)��iP��ą���!����N8F�l��KR��L�Ͻ��d���skw��1Q�k��9f�}���f(�U���hwNuY�|�EQ�$p;��(�F�2'�l]�e����Bqb��垍Ti3���I��ŊA��s��!�\��Kj�O5Y`i�g����Z�"�͍��	Y���Z� �hyiwj��5�9u����[Ma'�--�|j����w��T���3l��e	�q�>�{#��u�Q�wg�����_9AA:���=�Q���iTfI/&Z�_��f�Ə\I@�0�ש��O.��h��~m�b$խ>+!�D
��$e;�ѬC���O=�a�����)����4�P-� b����xb������@2T�$p���r�B[���-u��!c]4��,{�Y}9�Umо��.�&h�M�Uw&�"�0L�ɘI��J3MrW�3�)�S�����X���\*8�� ��xkX�(�� �Ma�l~���IaaIR&�Yl���acn
B�B�y
�֪&�0)'Җ%Z=�ET=�Q�y7�>��L	��()���.�A*Y��څJL�'x�8p���T�)���ݮ�:'Az7��>�#��ɫR�e4�O'nV���;k`;,�o���r���)Kw̧l[ml��gT��^�q̲pT`�)��!���NJ	�B�*�ZC�e]q�֜�T�*���� �M�R�l�zH/�m�BN��q]�rJ�����`��@��u�1�����JN����X}']ᒀQ��\���^Y7،6��Rw����ǰ0Y%���I$R>x4M����$I�c	t5=� ��M�2a	X3�]����G����Kt���Z�8E� H�k,�m{I��[��FY� �� ��� @�
�@��V���rG��y��@w���u!�$�����#xT�?��Ђ.� -�G.�km�A�(OPx�����xN 0@HB���G��hL�<��;�� 3�::�DQ�G�:��P��U6��1��:B�;m>Xu�*(�4z�%9H�=/`�;��{���PG��:��Ԁ+ਡ�@PP$UQ���Q�葬�QrS$�i7W���:��l{ ? vW�BÜݴ9�J �\�ԪaÜ6SD(�ٍ@�A��� ����e]&�/R��	�"��L�?�;�^�����'H$v4��*�vA휻�*����� �ly���PV�PZiW�(����4��E �0
� P��@�� 썒���U��PGh�E�B�4"#�Q�o��i)A�k5&��J���

�
+���C����EQ�rA�PA����Y �	�'%� 4��Ȅ� *�
,��#�#��
턙������b��PqE���Y(QU��J�+E /��PD�A�iT�>����3u "<�8>g�|��"jzO���ߊ5�����o2Ӿƫm��E�� �)J�q�x��*e�����!>'Fg��(
�xv�xP��B《�TB�w�D�T�6�P�� .H�9
�Ѐ-(�J
�m(���(�
�H +�6! ��AY	NN6�z[�z�E�^:�ήO[>}}�}��}l������$E֗�̠_���$_m�x��f�"Ą�U������J����>�����>���f_��Oj� >���1]~9f.iX@���y���=�*�;����$ ��H$���F�|�1H�d��W���8�K'�}�D�Ӯ���,/���P��F|�Ĥ�/_��S��O���60���V�MĽ�IA��O�	���XB�fl;4�����8$�Z<���x̽�A�\vc���B�irą\�r�f�OSC���̇;�}o����}^�C/���_)Ɖ=3��RK�$�y%��5�[��D����Ͼ�����)D
snڼQ�<�kk���,$��BYm�XA��XF��hQ�!�
�-��~#W�;[�P
��g����w��/�y:����ջK��ˉ��@@�X??CL�9ꗋ)"u��8��'ϫ�$����+-c�=�r1V;�N���z�=o�K�T`��x�bhXD� ����[�Ԍ�%*���p3=i|��#	*��d(C�@'�R����}��|�R3{`!��b���[޷h$W����S�B|�DR1D��: ��� G�DI,�|cb�Ѽ, ��0�֔�eP�Z,��D|�'A@O�J$�SL_k�<\�P���cQd�N��S;Roĸ�#�VfX[����(��2�[[фD��SX��2�-�����n׮�}�iw��Z�^B#�o��hA��������<��j5�����F���S�\c��K�
��j�QI�5a��K p,�TW�q��y���D�ֵe���1�!BR�m����!�Q�x4�G�$�[pU�h�L�S�s��\!�l��a�nE2-��(K"��V-e1����&<Dbx�LL�iNH@��2C��Y|7j�[���)+abRZ��n�Bڽ9�0]m����X�>y�z�
b����Q$��]�ta76��m^���~��!/�HCĚ�b��޴/���w�{3J&�����SJl�c�ϛĬQ �@V
��#	R��)����ϖ�a�A���հ���m����ItV���`�ÙٻK*D���V^(��@����ٛ�r@���Kc~P��x��MĖ�Ozg{���)9�`���h�����8�n˭�ӂ�oJ���`'��璷��V!�f��\OWλ�hO*U�%"�Qa>���)��>��Ef-����m��C��㥇RO�-F�"�Nx�H`���m96����p�������<�<ćU��!I��]{�����x<ilN�g�x��Gů�è@$=o�H�����
���|�k�W"��l���I����d�}�ذo����fb�� ��$���g��&�� �;�y!b����_��<�����Zu�Jp �8��)���}�4Y`S�OnG׾���0}n��'�%I�J��!��ق;y�q��B�ޖ�a*�r�f�{�5f'��M	���@l-�e:��5k�l^a��v%��! �"�	�Xq�䖫��B�1$�c@���9;ZP����2�f� iD����ޱ�Mp�LYN��Z�Bx��R���5��攷�>�!��}���l�FU���1�����S��x�#�,=�e��u=f) ���ckz� D$!3J�X_g���I<!A[P�<�+<^N������d�	������x<���Zӎ�d6�5�O�i��Un�mg�uF��1�M�x��G��( '��88��.�K*��u'��|![,;�g��<����&<@��y�PqDP���x�FP�>���<h,R$!������g�� ��l�9)�l��H1<|pc���a%"�(�E��`�q�K#e���uQ�����G(�L�N@&�  e,�i�HB_^g�G޻�γ���|FR���:�NN! �K9��h��W�wOX�O[� C��h�dB�����E�F0B� ����o�����oO$r�|��5�b�Ԅ����tބ��d��XфVX��3��B����+BD����P;�4�[��ϸ����c�HI�3��辟[,��)A|ڄ!	�i�͞���zeu���o��|�l�J�P�}]Еx�<J 4�N��Ce ��"v���	�B 0�@�ԟ- O1gƁ.p�V�W��'�M�gz��g�z��ԄI��8@�}�sՄ�5�H�������x#�B�}bL�T��ZR8����2Rʡ<�W#�|��N�|O)�I�������!��&���8*/s���ppD��͡�X�פ��&̐(��uRPj�)����̑2D��[ƍ���VO#�kz�CC���(�\��T�>|��
#
�KH������Q��.��Ѩ0� ͅ��3�P�G�v6��ck��^:n����Ӯ����s��H�	��!�J���@�YT�H�Õ�'ɕ���B�!A����o�����Dao�9�z�*��c��G��q��{�mo�Rv!2�7�F���6�xL��JV�UJU�e#�
`�EJ!�r(�����TJQ��

M���Mt���N0DW�vdBB7��?;��E�s\���?	�I~`���}]E�x���]@REY�c,�I����T��	H�N�hA$�/&�	�& �#�^Ԧ��$!H�d��'P�Y�z�5�F[XZ���{�T�һ7D���ǫ�}���IڇH��ρ�&�'6:y�n�
�ٜ����G,﵁-q����A�Y;`�ӐY��8�)��0�S��y�(~�#��^׽�x�G��ծ��DQE�b���0�1��ICBRQKC@Z�Sy]K��bp����B�۔	W���*�X�]FT���Z�ɏK_�W�5{:d/e�y*�_J��x����r޼�c�ޞf3�;�"+�_/;fBM����˳��TQY�h5���q�9FD����fF�E_:�n�;L'b@)D���	�8��a	�5)M�j�PTcDX���q�5��i�M�K#1G˸JAc&�1� UNTV�9}<�f�Dh��r�b�E�E�sd���-�Ŷ�`'6��\*��OhkRg2���6I&�b7,\�l:@�(�nI�ٮB3M�r}y��/�s@��:�܁DJBI�ș��J`d������{�Ԣ�$D�BO��E���J"��4�
;B)J;NL�iS*�(X�G%�(��٣|�e�k��X�E�%�x�H9n��� F�������"���IX&VA�g &�1i���}�������_���M���tz?��_i�����;�?x������!e�1ֿ�7�{~�L�f���ٰ������69(����}��Z#�!}��ş��� �N}����j_�~����t�7%��-~�����R��1U�$���(UL�YA���ǥʇ��k�G�r��5~*��^��On�<��+�{������
��V�/I�4�
����q�эx��ak�ܹb�sӑy�cd�;��{[m�v	#W��# A  _�-h�U�}���rZ��L9�&bZ'����w3���E�xf�� z4,��o�"�.�Q���Ա�g�A����Z}���σ ]k�`*�Ǿ�
�����֊��X%'�����*�����B:iH�	a?�:���T����n��#�4
˛��+�. g���֪������/���I�d�0�IMP����_���p���[����8Ǭ��]���	� ��D$I�*�5�Z*M��#2/��y�2;�i�cQA�0}[�b���e���-�ϗ����[��y6*�5r�5��DyJ��W74z�mkI��G��b|:���m�̢M{���{9x�ɲ���dH�����+޹�s3���~rE2�$fƽu�\��21��b(�}��O���O������P�W��G߀o�/�������~j��Wu����O)ȟ�:)��#�u�HRC��	A� ��Կ�:��N�ć�Ԋ�}���^��
���@-Q�KUD)kK���:z���_�AyI�t4��Q�}�|.�hY,�?�$�� ����ًpڝ�;VU�cw��#8�����?vZ0��?	x�Z�p䌦���/Ț���&(:l�w��d����']JPD�����zr���'��~!av��>�N(�X��;���'�"��H:Q�����w�J�e;4�`��������S^�	j݂��+�_��b�!�ѳ���E���b>�����ڊI��0��1a�}6�2���Y����� ���:��x��.��Y
1

��;��>_�V��\d��U�-^L��
��D������zG�9�]
}�����B,T�MYP����eSYv?���X�b��nѵK�~kV�.�-��A͖�8o�,��ܗ0ǻ{��H85E&�!�=��IG�z�bIos>0�"��Qg��H�/m�;����M6K�S��Q�U��.��X��l<b��A�rl��j�����W����������3�8��k'n3�|���q�z�u���o❪厮r�3����V�u�o�B�K�<�k�B/��f�p�搂����AIP�_}����\��KYp��>	?�F��WZ%��ú�1	=gj��ew�f�	-}31��w��Ҧ�~���sb����= ����)�L�o�����/k&�W���R��5���J�,
�mᴍZ�g��G�1��q����H��&}m��C��s�79w)�C�ɻF��'.��bX(���rBidEOh�2y��6J����F$f�����aS}��t3)������i�ۂ��я���l�>�/��GG�v�c�1_���&.�l�\W}ܰ�~�
ݷ�)!BV*�C_�����w`ļ>�#oM���[-������5v�*(,8���.����
�<���~gM��V�*RAV�����x���+ڍ.��&-/���x2akG�t)oJ�;8Y���SK����c�{̠��Sأ��fR$���:n�q����a��^�v�7�-�\�)�����E��Nħ�D+'O�-/d�&�i�S��B]�� �{T�as�y��Nt'h��f�,�L��ތj�F,�80ب���_B��/q=e͠��C��,�'�w�lFkΖ�^&e�&e��%a�M}B�����~�#!�m3�wR��F���������:Z����Qy
S}�UFS����F�Γw�!������Ah���ҳ�U�Z[dR�P�L���h�@�T*j��"g�7�jT��9��m~v���
�!�,�^G��᷼UߴI�ފ����(��\Vk���v\�N9��_;�7^��>���=<J�4�]�k�,��M�`���,UT�-G�**ë��[8�Iȳ�{�,�R�(����|/��Xp�U��K��Ê-E*]R��sXq���*x��s\�[�5���@#��lsb���Q|�6�JrZ��Lһ��|��Ti.;A�x��R¶��i��X�]�S����ߔjl����.��e�^$vbL�P����5iH�Jg-�M+�ҝ���R�N$�+��g}7��}����RЅRD�(z��� �����Pz���C#7��Ֆ�G��b�~��L1���%���^{|<𐑮p�"O]�H1��@��u�����W�J$�[ ���`M&e��m	�҅S��E���ZJ{ R�`T�W@�ë��o1n봅�DQf�4�5wv��Y�L�.�a&)"�'չA��o��x��{oF2�-=v�k����8I�� R<!�J=�^��}^�76O{r٣�ݔ�|��4�}{��(؆
=+�<7%�E\��cS��dJ�E�4�4�H%O"L[^_��ܯdI{�|�y�L	˚$�I���<q4wp(���wv0E$4�^�R����ۡ�d�IF-�&��h�������\���۠S��{;<y�p
�#��e�v�fH0ɷϹ���0a����d��-��/K\9g���zoNAF-}�/K����rR�%'(L�L6�����o]{&Lē�t&� �{�LL��v
J�����.��W	+��k�o������~�ou˳�|~�:~������{^��`��o�|5�>˟g��]�B�O�\��v;h������4���*�����2ܛ�~�E��?��?��(/�QeR���?��x~�����n���3ϛ���C$��K���= ��(}۞w����A�. �]����ـXcw��|�3�\Rڤ�����s�5�PB���x�3mog��
@G�Є�<	v��"��(�*��a9N��Xg�tr�s��X�5E��/3f(������a<��A��t<�7�*K��y>iY�"C�`8ŉr.p�$L)p�3t@��.�ɆnI%���rxpv�Ɵ
��y k-4���V�A���M��_}�Jp�-���\[ �Q�.|IE�jz�:^1�(fa�Ϩ\�2�
�(Sz"�wl�]4�$<c0����΀x���o��*���K�l�J��&�(4+s0��L�X4V*NM �F�,kf�=9Ď\B��[��l����ɔ�MaQEB�����B��7G�9��$�k�=��^o[���sU.,	�<��Q@�S�����YH�Q�EK� ��`��L��d��АÀllKE�W\S��+�/���hg��%�XK_4nC�E���Ĉ��÷x��P^�D��7�a�a�.s�
���
k�'�-�mQzu�S�N�	'8����"�$� @�����ǌ5.�f}-v|���d�+�`g����ME�H�H�J5e*sb�o���	��;��Pm�c*�q]���
�/+��SE�ѰY\��.�T�a�4`K��qy�qe�J�MH��
s��8�/XC;r�q�% (����0]´��Rk��8�@u���$�j�A��9�lk�R���7\2tD�h$�� �Ŕ�f6I1��d@�(Z�$Y���U��)�(� ���T���r���lX4��f�-��~�˱��c3���J��V��r��*�3aX�vҌm�/P�! �t���_=��*Pq��1E
z`1�呅�1Gf��l$���.�Y�2*�&"I�F��/00Z"6jm��&�``�l�ss� �h�7���z���,��"��<�Ç-Sj$�̲��:y�г7OY �����j����Ȓ�9�t�$tod�ƥ���
L�P�5�9"�]�E�U��Ϟ�czqO,�J�g�ǩFH�ܦ��n�V�1]��#��#ꭜ�[�����`2�X��U�I�  � aah0V#cE|܋oT�.w���}��]z������L�!cs]?,t��3��4bm���k�p�o��UmJP��@u+�P�����5��K����FE��qvFy�XH�b<|;�,B�	1����m��bK$lZf�������E��F��st7^ǧ�T/�t)����O�\RCRK�+��d�s���h�Lj�ܡ�� �����!� �L�����˚ǅQMF(o�th��	�kr�M2ROr�/wuwuT��f�)Q�^�cG1�7GWST\ݹ�]�$��A�K*��R�X�G �<����a�4����%K�������r��݌��q�/F���zsi�W-�vѨ&���
�r�E5ttuhն,$|�������b\��U�W6#V&Z6M�H9N�u(�'�����Ð`RE "(�DF��+�MA���-˜�捃m����|<��	��n�J��h��)Z���<��B���h>.j�'/���4[F��`�������쌘�PWӺ7{�o��ŵ�-Wë��	jk�]4Q�4X֍�'u]�Px�a�BR�%L�v�ͭ�4%m��s񈟉P҅�`��lcQ���cj"�����Am���inlI�v��wv��',E"� ps��+��$�d�NR"�$NI"v�tt.K��]�b���ss���k��]�6���8��"H(��;�+���\�E��sE��[����3ciLd�&"����'(>�Q��8JH>d&�s�6��sni+FI�����Uʼ\��vܭ�h�h*}�k��)��K�;½��;��M��"�+��s�T�(��q8�P�1��f��7�T)AT���	I޹v���^1`(*�k�c'���-՘-)H�*t]���&���cb׿��i�$��
��>�76{W�Z*"���sx�,F���b+F����|���[k���P�]ս���]Z:�v�Z
S�Jq���v�L�D&Ё����ǎ2���FE����6�[��sE�4	WR���y�˱���d��h�&� -_��ER�H�*R� 5(PuHơ������c�KE��|��=v�ί��!��U�M�X�W٫r������\8�%D�TD\���Ž�(M|��[�s�6�QcF�ԕˑS���cxCyQh����`x�81{�|]=wDO�pܹ�����]0�dTVM>��od�c5�6�1m��&I\`L�D�rEN@Н��o7ú'Ӯ�2z�Xؒ���>�����j�{y�$%7�sQ������h�����F�e��DY�<�o�\��6�<MAQ�E&�w��`���ޮ���ԑ�2���ڥ��j�CR&HP��$5���&�]�m�U�۽��0bƒ������O;q�E�i'���Ok��sXط�񷈁mb�%Hs�eJ��9J=����)��@��ч4��Ar���h�,D��&W���ٷL^�h�4�/��Q_�^-�}��d�:�(^9"P(t��^�lNR�� QxF�{�Pv'J4mo�r#0� ��:�E^�nj,z<өiWy��#�$�WRtI��lQ7�D����ExB4��`yA���<.hu؅k��F�0Ti���ծ�/^|��^ ��ۓ4��'���Q�-�X�Rd"d	�)D+�U�����]�_k��W�x�7�7��b�R�ܼ��6!&�����FJ$J�]�C�e�G�6��>�(
���S$r$L���
��S�P�w�E%#CVc�sp��LT�����Cllh"a������M�rM��Q5����^��W�;HP5�\����;B��
�n!�U�z`sX�:*"M^��A+Ӑl�܈>��ܫ��fD�w#3�� e���뤯r�!�	A�^� �&�F�C��䨝P�&��ט"j�nAU�/{�{uҢ�x�c}W���D;�hN|�׊�o����^���8&a11>��Μu@jL8fs�dJ�,��� �E�iy�C�D�]B���`\w�Jd�IF�'���UJQ[zV�W���$�7�((��%�6юfg��	�:�/���=u�M��ed��ۚ�ʹ�kd���w�yA�2�@��MB����.t��uA����x��r���lQ��^O��M���"���)
K&��W.��	��r��]_f�.�a�� �&A����Ԏ�b�^�Z ��T��08��)\�!.H�{ܠ���#EW��Xd��Q)�q4Ƚ�d&	=.�GR9�y�W��\�R����h�(o d��u R��]���d���
��z,�Q�p�����H���H�� gt�[�܍���b��p�}���7��cEr�,BZ/N���1+��"�k��
�X���@Ĉji@��S��I��hB�"��iu�A�-w˭�Q����r����.�������y��7y�#!�G����z��@ Wۮ�a�%{�p�ܫ��B��
G%S��
9������A��.��'��0mx��U�k��WkAh����_7��Q=�sY���H�N��c%���н7(G�n2����e�ԇ��e!) f!6�j�<֠���R:��5(\�Ю@�@;�r�@� »�_6��4
\ؙZ�>��v�`��3�s���Xư�0�ey��ˀ�}a+K$�D�.�W�쒾�u%���j����ߌ�$������>2�**�<g�ʱ��}q� �E4D194����8	̨� �"�6V��Ƀd,J$T��-�_�o�i��?(x������������=hwd�'���{�}璃�|��O���v>,���Y��?���8=?��,�O���{>@_y�G/A�N'>fkZ;DsE��r��/:�6v$5 v���|�M��P�8թ�xp�Ԝ&��G������@�6�~��~���O������w����?�������@w�� g��=�W,R?��������;��~�a.���1R&y����x�E~�?������I��g�I��"��K��Y��;2������h�!� ��/��Ϛ���h�!�lxۯ"���I�e=�J����;C�$v���7B b�$%�!X{.xeh�D�:R�m��(O��(�-Gz�R�ٰ�b��)�ٺo���x�7_w������O_^�f|϶��-�}�w3�F3��b�xE�~W!��U��g��,l����\�e���wI�%A�W��oL�^�Yf:K~,�/L��߫����m�zN\mx_S��vɒ��ebYl��'`0�(+�7�Q4�߼�3��S ��2\-z����j�׶�Y/�
"��.ܲ@#0���-�D�C:z�L��6�uBv�Q�x'�����|.�����aN��Yzx;K�f��F��j������b��'^���[����F�c����'g�CI�8�WǄ�����x��(�rո��3�����P0z�������Cg8Ҟr*��E]+#+���d�Vb湸�n��uw�iȈ`�����}/�>NB��x�Z#�����@����KU�4�LF�BѸ�ǽۢ'}�����VPg��n9$�Ƚ�KX�,��
���f 48>��/W���*���^��a�+���0F�B�9�1|jx*�j�>�̑%K�M��%�>�а'F�)܏�>��g����K�L�g�>�y�^ѩ���\U�yG�i��9Sݶ�٥f)��E�C9X߶���cH�Y�H�, ��V�%�9��{��y��Yr����x[���wU�nu8�ı�K��I)W�|$r+p���^ý�bh��]�Da"06�����v4E����U^�3�:���ך�'�:X!eĈW$2�´Es�*5�߫]F\�K�������<Q�^{jr�������S%R�	�֙)0t��I� �9?~t���遴�|�_�)��|�����!�{ھ����h��QD�@�e^ف�G��4�\��D�6t����!P�'��^a�E	����څ�^&�W�������5C�]@��Iz�>|6�y�]������\h��z���]#,����9�	�}⪙��FK��f,�0a[#6{3�U.��P�5��|Kj��[��25�Z���a�pǒbJ)�����0������lr��Bwz�2�|-7�'_p�Yp=�d�v���á�$)%hϖ&gOZm�-����pD���jd6�ӌ�q�#���Cx��}�Q�vFo;��Mw��a-���,�_\����;V�a��P%�� ��{�ܺ±�l�/~������b�%ڪb2̓(uU�Ta
9b���	e��`�n�}r;@��b��֞d�۹��푶έ�ϭ������W]a5�������3��=�j�ge�	Eʁ�X�I���)��<_M.��>7�k�d�A�3(�7|�,�H'x1R]eh���-i7x$���3;{I�,�~���Ԗ��~@���Pm�c<���9�i��o� �""�"�
��&t/2W�`�@� ��a�~��z��|.��&G�vU��3qېb'w�n��=]��^(gC9�3��~Z�=eԛ�I{s���}�x��j��Pu1�e Wz��	��5�xU��<2\#��ޣac�*gҧ9���S�L�ӷ��zzÃF8���v��Oq�.��LC��[�k��8��g��>:;�o�!�ߠ�*"l�$�3���IZ����e��ɸ#D��oJ��KC��ĝ��~9�g�9zN�§F@��=��+@axq��#7�:�?s�c/'�KI���(A��v�LJÌ�	��\>:���1<�q+Apn�뫽�q�=P��$#C��c��c޽��?G�����>�@�����+�+�I �O���� 䉧�������%��
}�����Y�k�����dq�|��q����� 7�������?����t΍0�������$��(��FD�����-+a��X�[l3Q��
��>Q�8̉m�/+��B�R��|�Jr��|Ƀ2��"2�2�ݖ_3H���00�d�i4�;��2��E�	�	p��_zƆl� ��$����h�� ��j�:.��ihp�5���'�8���; �$�#�7�*� �wUg3��2�E ��8�6`lʚ�#-$�%.@��YOh�O��c"q�HX<SB�E0�̞��pAe�:� ��$(R��Y��)��Y�����:&�V[,�۞v˧�J)�:A�0�)�O��P�KІ�oOs�m�5�S���`,��0x�k21��h��r/D�c���� ��0բ�e��+Bo�G0�e�qj�*��\��l�[4��W�@W�f�( �W�`�n���*[L�G��Ҳ������$ХDz�<�2c����Ax�tCr�hכR����ɘc�HɔʳA��F��R��U�TL�����s�<	�WUt�hl�0�0U�87N�˶㪦::�bѠx����肤�Jp���UM�N@�+N���u���X6�|$`�)Z��"�A��,�fiV�+Mw�p�A`�Q���lhVbKZ*�2����%���9$�6 �xu����V�oa�l�b���P)(���@�cUύ�T���`fuq����[i�`8�.����{c�����]� �d���n$���1މǋV&��.-z��lpz��4�-f
W*]��q[�	�
d��P4�����oB��fF
.r����1�EX��=0�}X�pcmB�dh�E��'E}̭zj	x���0�L�c3�S4�1iP"�Ly���;UIf�*#5BD!U1��-��N��. fg��$Im����(F�0sWd�r��IzL>EE|��VR@�]1��͍h�\X�X��s%����0A��n{��x�����I�Q��p�}��M��5�7�c�<K~2��)����6���NЧvzQ�y�(��S�� [9���2��l��Z�ʇ��=_�~�~���k��/���;_����m;�7�\��B��_������o��,V�������?�� ;���H�w@�A�C��ΛmlI�law=�x4P�5HЗ��5�J+��;��R�V�=?���;���m�Q�����gj�AxBDEAڮ���k��b�J�d����v�Oy&N��olІlb�9m��АC���@xN��w#h�gP�����B���is0�@� Q�^��w�g��/���G��/�����_�7�@��_��?����}s����1Ɏ������3�c���?����>�ڶ�&����]���J��te���f?��B�E�������Qe�q_�  ���?�(�ُ�DX�~���wYS��ῷ����G�
w��-�Ǣ:���DW��]�/b�vָ�`f)h��K�J"8���md���h���뵲�B%�|��ڑ+S@S�_ǉ#��>�_��#�	������F����������m�l�g�fW(h����q6��	h���ƃ�+9~� �6���lƩ�=y:��?#N�K7�E�?^�{y6"%�@�x�6�;*�c+�M�F`yk:ؐ�@[�V��gK�z<x0*t��>aUp�|����2Pc��n=�NW���Yu�heW���P�ZC�:=Y�lY<,��UK�":���Eo`A�����c{�]D�'1R^����;^2
R��u� 4n��UO�-b=�ɠ9D�4J���v#c^a3}ZqHy�im#�=���a6g�)�QU�!����沠�AB顠��W�d���aCƿ���y�	�O�0S믅���`Um����z�8�T�,�gJ&Vߴ�fٛ���Zj�
 ���ʂ3�%�����#6>Y�!Q��Gv��6V�ף���xOFP��
OC6�ʡo�����ݗ����"��7_�^���='��$�r�{���e�]�Hu�[s	(��lJ��+p4��?#�'/��X[S��Y˧��>���a<�"�'�!����s/����m'o�}�PxmJ6��։Y�M���i�k�󞖽���`�z7��ꪶ�b]�z�&�(�U�|yQCϭ�=-��\�%h��6�{Jq����"wƶT�T�v����ȟ�Y�?|��@</����t�ՙc�7��`��ݚ���d;�ݞ03-�/mq�Rv,]④Kr<�!���J�V�`h\��?/)�c�i|�/E��N�t~�9��H'��x�}~�i� �~��(NZ+~[p��y(�=+�	_3.�p��~�\�*���I��蠻 �~px�@Q|���6kE�~W�
X9�K?v؁���V�;��"�]��\{xq��D���h�E���D��$״� i���"x�|����3?Q�r�Kx ׺�x����wU���0�g$pRz>LO��Hq���Ƀc-�G�' �{��M�_�4�dE�;�5��1 oĒ*�ƾl�ly���������0���n��OYJ�GN����+���M��-ny��mս�.�ǀ�ͣ�B�}��(+Sב�M�{O|���?em�/���w��ZŞ�3`����>IP�,;� Lýz-�U���N4�������T@�)�E!Gg��е����}��AH(CB�)#������Ť
�Bff&n���*�гr4�8�Q��`��Wpɉ�T���J \"�5C���@��U���W�}k��m*2?ae(�w�ҰuR���+�iG���Q�[���%+���Ȋl="�-\cO7��"��S�����/�/��>ԎdN����k�7�q1$��W����P�M1�J_kE�!~�1��4(l�'�O�GnT�ų3�J�ϗB.\������[��h� S�;@5��_8�2�cW-F�ɶ����7ag,է�>~�����갃C����=��')Q270�G�2+q}����`�ߦ9]h���ݰ��ǢU����X�����l�P���:\�#6L�B2:�`��贸:
U�Q��U�B�=G��Q<[���&a��
<�3��AWw�R�K��D��mj3�;�A!�RC:�)�M{�Puab먥����:Ϙ.ew�߷��O��a^R�~.�}��Ű�[,�5�<��(\n��y.�����DAj){�}a�� �u�XZ�M�UX�3i恪-�x#s2��ti������)�/>S�2�gw`^�*�If4�d�C���+*J�/R���MOy�Xh'�����z]��al�Z�� ���������Su=��>Ȟ��#@/���e~�_(�~t /���H�~�f�8b~'� O��/���:B��\�o��H`���;�q�X�7�~ԱO����iB	�� ����0����
2�]_�tD�,?�P��(T�O���B�,Or�IN�zZ1 x�2����94��D#zH�XD�:�_)�)ID�-Mu�H�!���H�=�p: a�B�}�ȉc�PO�Ǧt�Xx~��E3S�U�0h��fO��� �aBS�a�iVN�`F1���@Dnt],�[�F�`J�$�T ��� lWR8�����I�$��r,�"�ք� �TF���a��i���~q��d�%�VW1�D����+Ca�"�A�(��Y���2ŀFT�XWL�R"FTh��H��q�>K�/�����Υ֡�FX5��"�	'�v�f���(�Ӎ�	T�t"��踵@�Kd��rj¤���.�� �Vb��X�
�#�4/^�����
�z��	Ɉ(�����x�Q�L��6�N��
�pę�ΒWH���</�D��"gB�%a�d#�����3(8ό���8^K�eY�XL l�95�@��=�&��,��\*�B�!�U<�������R5F� �D��XSih�9Q
�p�֋�$PE)�,H�Z�|q�4�8z��,�TB�(��H�C���h�<m�.&�u�\��������0�5}��:ቀ�sZ�Z̄iYe"5c �'�
?�0�L٫��Bv��i�+'Z�挂�$�����(N4%
�E�) \�2��`�w�r��)H�ʛ{c1ShUӲ���a�Y �U%%�Ic�����) ;"s�"ҧ�a�XkYCύ$��ÅL"�q�#�Y����}H�|,E[�4x�ğt�#=�M5���F�Ҍ0�L�9W�ǘ� 0���y6�&="����dJ��XLR���u�� J- ��- �lוl��-��|�"<b�@�''��4D���kV��
J<�Ȯ���g}!��?-�*�*���C��,��6"fv�ׄ5�rnQt9c,`qT�;"q�`Q�Z�,�|� � |Oo�>t�p�a��3"�|�3O� . �Q��LR�0/õ�*"����o5kV�<K��
<��}_�mվ��@���&#�E�*P���r'P
�4
���s��o	� ��"?A'�B��;J��)��,�A�hiECbUSS�(�u*��o�J��U��6J��s ʢH� ,���#��_���u߶_����~����Pl����~��[}Q� �s��R�W�N��}�_��~D�%�~������F��}#�a��~��R{����K��>���M"��ܗ�-�0 ߀  �� ����5a}O͛�:2�\L����_���*�����"|�K����t`�&.{��-&��ś�\O/C6��F�ߡ�{$��^�@����ލp����-0�TT-���g�c�M��I�A�\�Q%�&6��T�X��-��=  �����������!�T4x��3Zo��� LA�<kw�^=xC[�Re� ����}�6������z"?����x�&����X�Ў(�M>��.�i�eXK����UT/��F]�i�'U�|����BU��ў�B�����/�[>7^�aC�ͭo������<�f���4���<(��%��眜
<��t��ac��\`є���K�qa�;�q4�'���D��V��cu����~�S�}�x�Wd�������ԋ��'rޕ"�
�A���c��?eO���<�oy�$B�VF�d5��z�v: �Ԋ�1�wG�4\�-tu�v���8�׏�i��F��;@���抑%�Y�'H�v�]�q$(�c�9J�܉m���=�cP�0^�Cos��|�,=���r*rYh9��<=�Q����݃��k-�z�T�8�33ǜ[B'W�8׿Єj�ŝ�p���������XWQ�l��t�;B�g-�ǌλ!�|)MNv�b1��Y�=��/^}"�I����~��o*�7#n� �$�w��4�Ru�|�:e*Pʻ���b;/�R��'����*P���֕Q\��?������C|�_gG�Q#�b}������g��s�A���v׎�YAL:��Hw�{<�"�A����+��H+�T��0^���Gd�������i�N�>��8�3���)Iק�x�A6�K$��G�������Xy.{y(u��umM����c�8�H)���m��"_&�{�>Y)u�(}�ȕ&ɗ	ĔR�qޠ�:�ـ�*�O}�ɳ��A���.�؈�$�ET#���JK�,8�i_�;�l��>�9F�Z��;U/��R��Qw�K���;����lPL�����֏�;�K�oMOB�lt'��\�F#8M�G5�9e���O�~/�G�r)��|�'�o�9�B�-F�i���`�:���I+��p����-CTU��z�RS(��W8�8�rR�l�>ff�J�wQ~�G�h�lZ^��iQ�={��t���t��=̡��H��N���1F�[׉m�r��q[2��ʑ�� L��!Q�%Z!^�q-S�u��lZ��#G�:u<yĄK�*fX�Y&gZh��X������6�N��N���EqAV�Ua��9�!<3�9Y�<�E�O#ߧkB��ԑ9�mc���sI���O���8�rbH��K�����ψ_D���=���x^^����c,/[�D����
����,�E]xa�U�=��00���c�z��(��j�`��k�y�k2,l��۬��55�rBf��������R�?��쓄t�N,���Y���X���,k޼�Cf�Ly��G�	�d��f��l�q�!k܋��{v��8/t����K��w���'x\�]��镆s�>G0�':.5
��s{��č`��)egs;�I�CGC�)>7�*߳h�*�L���dc��몼�z�;��7�T�xo.A!;���y >=�J;�&��_F�֫3�ͳ��[`{Z�]�x[�Ci�	�g�>;n��цA�n�̯���~%�x��q&%��GV�0Aׄۧ�u1���l�e0����ç��u����I���{���X��,8W�i�#��҄�h�U&g;l���;D�����1���n���E�J�,'퇡�;��.�}L�u����"�[�B�Mf�p?E�7�]-$g�}����A��r���%EW5V[�;��Z]RA�Q4nrI�b����R `XFE)�z��~�����潯�|�o���a�
A$�����7�_��iM�K����<�G1&�a���@D}&Q�D%}/���|ϩ1��!a������A"�>�/4"�vw�:3&�Q�(�iq�B��@��
�<���zˤt��E��C��Tb��V�F��8�A+F�K��Ȗ1C�R��Ф��(@��CI>��~	�[�|q�x)2�iGM�0X�CEt�=	��W.�A�LL:���iV�~il�Zh�4	��b�/�LDi�ʶ@P��4Ƨxb�"ȠH��BaM,9�������N������)�A��i(�ې�Lh��W�Y��)�9
��dCaO."I��-R�L��S(0�! �(�%@�VC�d���ج4�1�6�5�ba�L~�_z( g�X7"u��B������M��U��(��y�-��8����� iC��6�\l���+��&�x6�CTh��� i�E(� 
	P��kB9d��b��FXr�[��#Y[
 �(*m�S]���Ïe�z֎A��SL�Mf1*�LtՄm�\�E��� ��
�b#(�.q��	@1V�1k���*��)y�Y����*:ʩA�wB0$��z�-�C,ѝ���((����]����LK�?p#P�U�[#�۝z*-4�,����H�( �Pd-��F`B9�53�L��T$�pG]B(��1��e�Xhq) �A��Db����iЍ�ǯ�X9d��q�7�,:���8z,���y�Z��)��kw���_j�>�
�;�
�&��6_�+�<wXDa'U�By��d�D$����(�#E~��2((`� ���Mgx����e%5f�RE�]��Y�H� W�S��f^=Um.JB���*�0T��@� n�"����I�m�ȡ��Qx�&I9�Q�=��sw����.�����]a��Ts=G���Q����[;Ey*�P�A�4�����	�?;����럯�FG\f�(�3m�����74m��� �����_�W���;��^��~O]�^��z��4M�o�KB?��'�l��O�@��>�騤j��Ί�
</�� ��A�4Ig�qf����X>��|��-gX�w�8����������%xZ�R��`�������?��M����b����CP�W�b�>��*��#f������[���]�R��㬣�gh�s:���v@̚�^,U¨w؁�ֈm�m�ߕ��/%ͫ�ʯf�ד�������%)p~
5��.^�!xݾ�3K����� %�=1�q :О�̜�����X_Q���9y�G����3*)�H�_g�����7'T$O'�ޕ��%|�b68t!I3��H�1+�)RV��ZA�D	)I�8.�ʘy��o�azQ�
醾T�t�L��շ��iY��fl�T�~t���k��2�F�d�P������9���<���رr�&)�7���3�n���b���mv�q�7ب������;�U��4��9��P�}�nՍ�PF�OrL���+���x���k̀n�'��T�0�r���B�{�Gf�݃�?�FN�u���S/�Br��Wi/ԫ�%��Թ]�l�|�����@'{aW�8KQ�fK%�=�Kمo8���Յ����aE���dy���jL�����y����_i��l��MTU\Zi���
���=�6e	�����,�½K����J%� ���T���`^7yǁ�T{�� ��ҫ���� �lL��e#)392���]j�}�~�#]�lc~�܌
{Abr�N=ϠV���C��e�_zZ2��B�asT(a�5W�طv�.ZW��#QCՄ�')Lǈ�;.Y~Kv7�#�ʲ��ǳ���U�o����.��
Ś�k�LUKS3a���#Ĳ��MG?m�Z��(;�)j)!��s�˨��n�;��|M&��0�]���7�tϳ��$�c��ϐÎ�1���?���X����b�b�4�S��,"��&xh�'4�̷�.��Bx�l��/^�TY���	���n2g`rlmE�-�t�R��ۓ՘��&��U�<��ʽ��Y��&�L����k����IR^Rg+;�0@�֓��9=��\�V��G���Q�e��E���$=�/��:�iB��6���]WP���8s��@��@弿l{���3LC,&�����2w�'r|�δ�s��9�^�,��d	���[��YH�8���.��B�|+�<�i��ޗ��9��Dz�"'ݗU�	ܠ˅m�Ip��8����9���՜�d��;�bw���`��U�S�
��>�gX��y�h��m�^N�/������93��}X���ƣ�S(l	j7�+�؆���~�a$z�(���^��7C~�'���U���W�D.j�џ,�7�<� ��.PsyL/-����L|mR��ꞵ&k����Z�y`���ޓ�jnӫ�AK�6���bʛBr��w<M�6>��a�]���1M��vD�3�驮�Z���$���S<�d��ܰc�A��,�J�8��&��l�RtDXq�2gb�ǰ�V�M\ju$��KK��y<\�8UE�X���x��!קϣ�uh�p�s_d�2�c�U'Y0�l��F�Q�K�^gm��W���$��g4��{~n{�Z������+��Y��yn�_6ʒ[(w����l��uw�9�ITN����E�t'6I.n^�����`��\��㼭$����(�f*q�������7��9�����!�*tϣN�	�1!h=�&r�Bw���̨Y)�(:�ԉ"?s���vz�)v���2|)e��Т��Γcf����iO��!l�'�������&Ȍ��v-�MFN�d�o'1��N��V(�:{ЪxSiE��_��"�5�����y;4c�J��>O������ �������7����w�#�͛��'���䁾���W�0!F�E���&}�qD��|���?L�4p���������,�`����VO�8nɮF�M2@p�OL���"��yH�䩀5@�De��i�4��P<�h}����r^d��EM�Ӛ�Ť,TS���fcIX֫� F!�Y�*�IbL�]��_1�*e�1��K�'Ki��B��J�3c�!
2�!]!�Q�RJ�<*:�!�L��<*�%ܝċ4�>��\R�5KNr�U���!T��t8A��>�#P� Z ��v[i��f��E`�q�a��RQ�:��1�huPTQULD��D�t8_9�\�3�f�R�D���D�1P8d���)8� g�	J���˅��q�W�"%2�wZQz E�f�ٌQ�x�l3�Q�D���Ω�H�WЉ)�(��� e�h�:RD(��5�:�J�"l� ��,� �	⚂s-f�xф��
Ԧ�Q���FhL��6w����8Cᤑ�T� ��p�*ܔ���q�`P�i%�2B��@J�"�Mn3Lu8�%�rm�@H ��Nd�_fT��66fEE9��y(��A����#�-�T砫馻P�MR[�)ԐqpBG)J��
2�d��2@��F��<�FS����-AP�DF�T�.)Hԙ�/�1�Yr�K�$�ȍ���3 ^�O�rc��"B&�X��i�P(�#pD�U�����[x$��J�Ue!J���3AU�p.�//n�F1	������S��=���W�o׏�����NG����c�x����y��)�Q%\����� �C� p@�t��"	��ٸ�a�0{_h{Z�gۛ�7��s�������������q������_�N����/��_w�y=���"(if�9��T����e��LV���n�du�f��v�5	�UI�of�����X�x�L]We���.���[�1�+3zݽ��#���T'�zr)��I&�f��:���3G{q1�@&�q��I۵
2�t%����
�/:��9���u��7�T4�NN0�C����uy]_.X=���.~���}��w�T/.�L�t�϶v���;��fO4�٘��Ks	�Z��;��t�p���	̏q�V�Gn��UUy[Z�:x
�ے��&��\��'��=�
r੹0�E���YkGUԋ��rhd���yV�c�}�tښ�W����4n�n�c"�h�F�!KMGUt���2r��LFc�s���^,��4�Z�k]��E�Fh�]�����a�8���Z�[�z���WR����/���W�TΕ�UK�3.�ȕZ�������&V&n�hj��[umS���8�.}69fww�pǧ4VF�vg6������fD���l�(��l��xv����-���d
��������w�)�M؄#e�J\�.�n�a�ztv=����(8�5��҅�V>��n^0��32�ͭQGJ�Ñ[[�f�l�s��l���'��S�9?�<o�"p��¼:��A��E�|�=�^��^�����������_���7��4��S��?������!�~X�;�-�	ߚ3T�I#��z�Q?�7�����t3U�]Jc�������-��)o�!�P�?/�o�}W�Hr�/�~�����[7G>��p���fc�Y�}�xԇ�2�n
k�Q=`Z�!�d����鮥/E'�2@u�J3�}BÎ�:8�'sΧ9P��"�P��k�x%X�B�e|v��YL�����J9y�hL7]�~dmBj���7�3�jO3��||��K��<!5�ٵ:�i���y��ES:��S@Ė�wS���>ŭ7|��$ݼ����p&Gw=g��,YbdqE=a~!���3g��`Z�0��C��[\�����I�h!���W�4�ka�$dz�z6�H��qڂ�_�}���j����nRn��nu�Wv<n�䒳�X�����/ܕ5����kyLJ�b`^S6�MY"i��2�*�e���~i�{�.f���mɐX^��Z�$��*V�!�[��c-���M����7�9�[[�������x-#�t��$�Z�����-b����M��Mjg�X��v�ϗ�`�I�mT�|����c��>EtI��Rɵ�	�Z��|�T���Hy�t�f h�
J<!J����FX��>�[���w�6�爐�iá���QL���M���+�|Ы���F��de�� X�����f9�Fz�LAba#Z��Ԅ�b7�"����k�$ z����bb���i�[X��nZ��B��Z���w)U]K�*n�xN�PLX���zVX*��_9�A��>XB}�ʒ��hmQG�}�ٖ������̱m��w��UF��p�@!������O;K��Q�e7{��3.��/��5�#��/�Oy{J�������a��to~U�n!�i��ܱyk�����o�ҝ���}���nu���ү>��vJgr�xނ�I�w;�O�ކ�y��O}�(��@��y�}[����%��{τcV�R�\��.!���m���4EA��M��/�φ�e�L\�yV�}�7)�h]ZG$U�?y�i�U��M^�����%B�Fc�gs�U���L�ى�y�6	|^�>ߑ����*@����9��q)hQ+��#k,���*� 9V�KSXX�n����9��e��ׯ4����g4o�������'ԏw:���E��C�<�7�ٷ���r�Ψ٬"�x�z𞲯ݩBN��a�Ac��?;�o�V���S�SM�E�i�SRWW��j���%�߰&�������w�
,�@��t���M�g�D�"h?�=�W�v��I; ۥF�RjWG�^�i/~2B������W�B�h"!e�/��R�b�,MWOG$:p��j3�*�x��S��q /��^��K=�"]��8�l{y�i����}�LY.����iu�>ypi�g��\A�#F��t`1��KQ6�xl���Cu��Q��)F������w{iAWm�����P�yw̃p��n-=v��N̗ |^�&βq� �F�&�{�;�#PV�܃P��޽���I��2F�& � ����[<E�a��^8�Q�=Ϝ8<f$E�	��<��ikYݝ1��$���;}��+�i�zqS�2N]+]�|����3�%� ���5X��5i��}��#�/�R�
0���aJlJ
�][����3�w��R��'�;����Y�>f,F!�����B�jF�Ou+o,��qw*[��ӧ/�2���~9w��W���y����.�g��r���ہ�}��ɶGݾ��G
�p�5���}znO٭5�O6]��0�F(�g�y��HkTʰ��C8׍;b�����b}!Jjz���э��Uk;,s��D�L��9�IY�s>��u��Q�����[�2�N��z������c|�U��X�cR1{/��e h��J��j:l�-�$�Wg�E�~#�b�N�77gk�'
���Drx��a
mj�J�ԯ�!�&^OQ�g�.'�>>��@�(�߁�>��>����Y�?~I�����gsJ+O���~��'�&G�?�2�O4rl:�$���N�(5�\qV�[��)8U���0����}�	J����W��Z{qOm����5���k���~�:��[�ի���M������ԯ�+2��sQ�G�~?H<T�9!$��R�11�V�%�ޕ�]j ��F��fYWf!�Rr�#�h�E2��Y<XH����o�C�9.�S-�N����<==~������Kv���m�1{�&o���T@hC��/4t�,���:�N�zW�ɠQ��W0T�\�S��[�Ll�5{�	۴]�������k�{>��o������ediS���2EcX�#I�)����yM��T�9��4�$j�F��RUm�7�A�.��M:1��!xǚ���l������~�dX��[o�|���~s�ׯ���cH��� �X�8M#�6�}�LR1�0M<��E^v�D�`C9(��ߏ�ׇ��;�?��Ќv���e�џ�������Y
�C�HHt��@�N��$|ЀCJy�a�� �ˋ#�}R�]j��'�4�,������_��}���|N�C�������z'�����C�q̿+�hy�v����~"��~�3�?���<�ã��W���~w���������?d���Xc�S{D%}��ν��t���8oS ��TG���~�v�7½}ݻ�J	����,ե����m��87ʝ 7F��,��u�x?����4�q?�G�*��IW�g���X��=���D�!|()�J(D�}j8 �]�1��(�?h��iH�]�4f)"QJJ1X��Etռ��+��s�uۃ*%�A�ݎ=,�f�@�U̮z�#�k�m_���k'p�,lu>�f^�<��`^+{����7Pi#�ft��<ie)G*B�C�����_3Y�5sN\�������r�۝��%lpV���l#9A襕1J,T��{n2hB���c6�	yɩV:*F�o028tn�D�ҩ��������'�A��,�Y�x���P�/\ �2���w�Fы�띄F�[��S�"'�."�.�wg6��qJ�\�3.���9�W`B6����f6o�_ v�򹩀y�Q��%��ދ�-��}���c"���ضS��]y;OJ��d����g=#y������BrLm�	3r�{��oF1Q��r6/����ד��#c�M��=L]x�Q㛗n�T��Ӟ*ҌXx1M�w���Y���wU�����)��:*�ޫ$�o�W�K�r�њ�y�FVc�ѳ���R&�U� -U���Y3{�7K�kw:/��{�ae,���gk���`�ǫ)tn��Ђ��^`�&-����WS��T[l���O=V�BΪS{[��������Ƿ���5ӭFn�WEj�X�;�p�x.���[vQ|�W/�N;d�gf��.D
!�uק��{������(�1�9��Vn�mT��zc$�ȳ��9ê��F,�VV���UP������a����S�8__T+dp��D��=�&ӛ髭��s�u��2c_n�3z)\��h1�.l[V�����:�2���F�%���I���̫��UWz
o-\��F��ØF�iۭB�L�
�'�>�@FՌ�#ΧF��5�q�\Κ�������,\���'��=�N�z�<;�[�#�sk텅V�ܞwr[�Uj%�?7=��[Yϯ}W��K����gyR����o�67֭�U��}� /�w=7�{?/��<k�=w��ߋ�?/���ܝ��3�����?x���?{�߄��<�S }��~�e�#���"�^ϟ��K��7�-O���� ���}d�bC1$��B��6/�s�vt2����U��2p���| �9xC�Y:�e�֛�q����uQ7f\�<��w3��l�����G�=wi�(���by��G����yE#��߫��Ǆ�3�D�.���=WY��nL�ڋ�N�wx���V��/�R&�&���H۹,Zq?(߫��rm*YI��������rŦ��.`�����֎x>� � R���<p-����8��|R��0���,<�V�	�3�H|�bb���r^���f�PH����I��sm�Ǣ�o^3�B����vZ����D�ܳ��b΃1D&�R�;�='�9�vd�ӔP���0����I��Hj�.�FN��'U���A|��v`e�<���Ԏ���÷�򍇠�q|�U%\;�e݅!�eE3����Č�5.J�U�0g���R�[��0뉕�4����U"�=v\�W����|n�9l�<�ggD`�����U�0����}V�]�/	�:��r�<�$�n�kd�5;�NX���[����X�Uل��{ո�:x��Y���OFY�2�J̋�8lh=�����h�k ,������Whi9ڙ�h&����I"(tix����?�����*�<�6\#@Q���xt�D�=�u�C��d���Q���K%1�j��S�g��D�ލa��Z}��wt���I�̨���`~$K���[�@����`礹��(�_;��&��2h�g����}[6�tSb�txI��!ݞ|��g�|6Дp��拲s�a�E	�8<�E�u��"T�>�A7��Q��Iv�&��V�V��+��?%\W �O>ِ=�I�7(8Wb������˳������h��	u4u�.�4W3r���i�l{X��vFq�^�Ge�k�(�ap�"�v�Ii���]����IX��,����h�E4��IP�L��N�m{�+
���0�1���}���-�ջF��1�x`���I|��zzz�'���&,%bð�t�n/�q�ѯ>눒e�-���]�L7(�p.���j��+��%���
x�b����٫��A�(���_t�y�m'���fH_��ie�&�%,�f>
�-=�($)�c�4z/��F�t���	��Y����s$#?�ť]�ʐ�f(s�u��+�e�Y�FAfݜ=�P��t:b��c���V0�FT�����O�!�/ڡ&�Y�5W2���-f=Z���A�C7IۃT��*!&�6FQN�3N��(�������x:9ڗ���2�{���ǈ��☥r��5�V)(X��Y����Y���]$�b�$!=�W�4vy�1�{ԧ�;���p��b��"����n�*�k#v5HJ�cW���׹@(Y�`6����Ϟ�n�T�F/�x}���.\,�D�^ȼA2J�,�	�9W��.��x�:�fKM���9H�iW����x�G�wW_"5m:
���2b�6xWk./w���˜� �U������z=��?2�)���^xq��<�B���E��%X���wKȤ�xv������9C1�ZA%Q-��ǖ�gya���eE�I�Ja3��40�0Έjz�'M�2"PC*:2Vy�c�X�y)��¡�N�6�:V��1O�-��)��bm�Lʦ�2v����I�H�R�\��Q4�t:B�	�Z �V547ɞ�qRdPq#�o`�p\���/��ux��7C2���A�;qq�%�㰉������e�>xV-z�wc�����v�`��m�[����{y\���,��	k�ذv/V��*�>�y=M��������O�U�M/q���T��3�pcj�DR�|�/�b؋D�=�������-�q�R���z�0ޮ��*	��Z�2,�*������J'�~�nJr�bq.��R�v��J�/��X���� � �|ߥ�����'��Q�/�~��Hb�7�_�����M3$��C؁4�cV��4����G�����0�� 1�hF�5�t��F� �Ih��	����.�ɌK�~������W�$q�:�4��_�8���o����
}&��o��o??�o⟎����߿>ֿC�l���iͽu=|J��A-��:8�68�Eh% �}e�9&!m՗Ze4��(�o{��w��,>��5��������7a����n�Oo�h��>��
���M�|h��C��Q�a��
�2�+����Y��O��_�Q_h�����#�z|F8-�^��O�M��~y�����s�un����ךF��[N2�����?Y�[�������?I�vo����N���e{���}��L�/�6���ߞ�ۆ�����+O����u����W���/�E<���{��ڒ�w����̐�����<��C+�>�w��	����`%�<7��v�����kG�>��7�q��>���-�������7;Cl��? �=�:��?��_z��c���m#*R���������o�v��,:�Ծ=��.���s��Y�����:�O^�����ߘ�������>���w�~iO^�QZ�x���+������������Ǯ
7�u��`=��b��=���Ѧ8W���K�N�)��;%{�׎��'��{`>z�NH��|��Oe��o�u�?���1yU-#JD9�?���W�z�8u�}�g�݌����=���M�3"b&��"\�����H�;7#�G0�����(�	!��3��~��e��9O��E}��,���/�������(����뾓���?�Q1ϝ"��oE�M+�����,A�B)��1�'����~��A`� >2�>&o�$����|�QB��mu����'�|'4��fM�qɀ�z��ms5�Y�Y�������M�%��ϡj�!���>˶E%�o��!4��\��#<�HH����{�����k�.�T8P���[bLP�#�{!y�����z����߸�N��	6���\Lvk���kM���{�� >   p��n��]�c5b�l<�b��%��,d�"�z�6bܟ.�x�'k�"��(఍iH���$��^��U���WE:6��6'�D�UCo�Wq�Y�D��z�1�oKڹf�H�S�0~�jQ����_q��1�d
lƎ�]�(�>~�p~�Y���S1�7=�J�ѣ��g��dD�K-Rb�w��쟭�n&�<��֭J!A����+��נ��Gl6 Ԟ�D.�¨�ݤ(�zͣ�2��Z�!�ﾻ� R�e6�kݞU���l
)P��d�a��
�t���I��VhH+���7zB!���J�����	�(f��� ���	q��C�ݏZr�B1��m��4��n�{F�I�����h2��2=%H�9�*15f�%���6��m��Xd4�~�uʺ�l��t�WA��ʊW�4��>i��d�%��c.+�g�������p��{�}纙�h��U<'��������ӧ�GC_3ơ�(�J/ߓC��~{�؊2��ƞ�,�y���hˊE��z�X����
L^V�j��΁��Yy���f�W��sd��YtR���Ғ/V�@X���Cf�C���_�s*�H2!�Qs��������oO ���%[z����]�>����8�Z*B�P�S�-��B�?�~��3}��x�QJHV&��̀jo:"v��M����l�8T:����iWDf�㤤y3�y0�7�T��W(|ЮRD«�ЅLchx��rOdt,m#z�c ��{�ެ���TC>�&G ME�2��?%���.�Y�����'��j|�j��WK{���A�Wx������M�����_�gu�5�؟��0�����QWX�\�8��|����D/�p�ŰmCA��+XY/�r�4�/�<����g�g��-��]��PƆAvT��,(�c|;!H�H��Ǯ1�ȶۓ�-�kp�zR�ۭ��6�oJF�	�.���I��aS��Ჴ5hCi����}x�0@���M����'c��l� y��K�;�b�[�#a��rD>>�o@�MS��ѥ*6�̉5D����9�����kA+�L��*m��Y�.���O]��)A<�wѢ ۼ�U���ž�zh�PN��Ȥ[H׃�f��S)�;<��^��K�m/.��i��3(Ps��;��`�[��In����T���Ÿ�c�Ue�S���������͋?�{s.U��tz
Q�Ζ�[(>7dv��}��4ْ����B��/p�V�g܏ �6��Z�Y8ls:2�H,���x<R����'�o}����|A0�꺰�[�`	eo�=������K&�GY:����y���}B��[(Mj.��;E9ny�.��)pa�]��rոp�<��~U�$|nT�y-p�d��^^�#X�e���)cv���!bY�.ok��.��T�d�I�=^��c�/xܜmN��zaFa�p���靅 D�1��'=O��p�k6;�z���<�1P(��Z�CR��.�0���KM#�Lt�Rnθټ0��x�ܦ_�*�V���i=p��:��M�Q�r�kY��M�E��!9�����\F�9 �P�i)��z$����#�����[>U$���,)�9�բ�? �w�ۅ<��WG�'e�H�La�fɇj��T8QO�����f<�N��4�ĥq� Wx0`ъ�$����f�ɸiUa��̶<X�eN��ZVi^~��I���Uu,��<�d[~BX�S�oʰ��"Ѵ�H˓�|k���x>���/���( ���J4 |~|�����7��ߒO����O��A^�?���䒘������C��QϤ�Du�L{b�z���-_lo�K��/�Xx^��}��-�$v���
Uxn��1����NH|I��Oz��S�~}�����R������G�5�խ��}�aoz��e�lz�����W�2ׄ��S��=������F�׿�1֯�������Z|a�����O�P~���]������Sh˘�o�І�{�U���|��:���h��k�:��]��u/��&z��^iO����j_��~O����M��Gc��1�B��v���Wou��r������_1��o9�sώ1���i�~Q8Og�|.{G�D�Ϻ=x�{��yk��!�\|ag_9���ǟ����i�A��P�s����{��x�aX�%����&��ݟ��)�u>��ח�s����^�ğ��g����G�o��>'L79�Xӡ�<�q�ɽ��,�������Qzڽ������ι�]cn��5�Kl��x|����;z��}�_O��tm�����j��\���Z���Ś�U�X\MJYQ��Pw	����.Ko*J^=�>��&�g���9����\�9��@e�~��/��x���n��_�{ΰ�	�z������>6�2�&��Č����ɶ�NSӊ��@���b�U�(�F*��ݽ�=y��)���i��˰.Wr7�I���ۙ�ޛ�D�8#'.��{.r6��#n���83��ة��r8�-�'o�+;���Lm�x.B��rv�':��N�1���YiӼ�j��Ŵ�5�����_S��E��ާ˶w�w��̨!UT���q&�#Q�8�˯6�ZJ�Vv�C/�!��<����=�u�.���,!`(��wK�2�����\ef���{5Upow�W�"�\�qFOKQ�i�7�wmV�x����gjo�:����ܙ��|�[C4�c��эw�:�$��`a���UPts��-2�������MqB��E�.���;K"Jc���s�nq��J�{;.\H�ք�sҵ��'-�������n�ˣ�Un�bb��XS۳F�N͙ɼ���Vj19U�K�ɺ6���R����r�a�RQ�j�:�M�ˌT���\�������������r�����]�d�%�iι��:gCh���r�L&5�4�r�B*���vX�w��(�Fi����,�����Ǭ�V�v�F��}�	�͚veD�%k3D_W��1n#tW:J&5��kY�W�rôj��E�����ᚵ0��Oj��5�t1B�Fq�r��uS�H�Hu0�^�
���/��=
��X�f�/�h�UkcrԜ����O.��uR����m\�T8;�ں�M�퉻�&�c�眪^n�m�EF+����s4��^�vl��c��vKO�O� ٧�r9	5�H�n�Gf��ynt��U.����u��`77��7y�i�\��u�uP��7��W�W{s�Zr��W�)�@���m>7x1P݇P(v�s|�����	���3�FPKo\�m��ðN��m�c:g��a
n;i���d�ή�6���2�!m7;+��TR�y�F�$��Uf��&�4(<F�S��C(M�K��v�;�,��gS{q�v]κU������yy�EM�@��S�"�l�Inj�,S�,��&bEf�S����4�� .��û�g<*Ri�a�����o{��1���9p\�ٰL���I��9�{���02�k��}WW�=&x?P�}��
��x?'s�>t�lJ��o���PMLv_r�67$�U��L^ec3�9m���S��TR��p�:[��\�!iUg#q#QzN��"�Q�v�Bk��S�2�T2&�GH�z��6ӈ���o+qV��4G�T���:�^QU���S�,<-�ՍJw@��5qV2��H���q�����܈!�2v�^����B�+-��*���&�+|�R2��DC�{�(�{9#��wݴ��ʣ��ыˌ���=�� �b�����������t���`ƮKF������7���c"U�G*e��v�f!�;Iˊ[k�51�]utRu�M�5�u _u@�Tw"V�`�3�]@ՂX�f_E��1��h��\�ev��s����VF�1f��Vl_;y��N�;#�;(d�yJ,h�m��nsR���������=y�4��X�k��f�;g��+�[��gGt �u$��3�0�dl�Vm`�"�P�dۉ�WS��*����VpV;�7�9S5�s�,\��q�`�9�:i�F�2n&��s���/�O_
	R͕YI�'��l���s��@�슜�_����kwz�d�:�]=�g��#o.�`�\�^dWE��X��)D�ʾ�:�*��V�6�鹸��M��\F]b{u^�pܝ�:#�Ը�zx�F��k��EaʂWV8��7�/\fV�]ʝ龷���|��9�5��g�$��t8��.��+c��9�L^�'f��u��k���Q�J�xX�V�K��ؕ}\N����J�.���Ma��ՙQ���3αVa1c���\t�\nЋQ�
6���VZv�MZ�F��0��1\�2�����C2y���r���1�(F@17X$e�f�mZ�q��1KK=up��T�N�<P������a�2)NI�����`+r�>Ef��dV�勣.��F��d�[��ٱ�/wr%W^�MNv��'�1iG��(���g!��V	���흚�s�[hÍ���[�w�Z�1���&�7�U�f�D�z6�N�\z���fu��1���ki���/�i=��9�<R�a �j]z��A�}�x�����pq� �9b�}۫4AF0��S<���:���X�S͌�v�����MwK�2��X��euR+�V�F2;#1Aj���R,ds��>d�C�	�����������$.d�n`��cw#f�R']C!��U�(�dN�fʥ=IJ�E��ۣ/���k������]�Y6�Xଋ��f���O���ж2&�Mu�f��f��m-#:�̹�{U�}[4:2f[��vu�7�ؐ�͋�x�u�;[�+3��X��ڹ�D�4�礊���.fs��[[�|�U�$������7*�FڻX�R�ˁ0Gd)Ӭp�؋�W�$f�'�ɂ�κ͝n�p8��Ø̜p˪�Zz';3�����ܽ��G�"9�ٟ�	�ޛ:��g,0Tr�3Л����m)���`u��{�U]��g�Ŗt�.���"=�/�0�����ķ;]6������V��Z��3�^���q��l���z���]di��HH9Tݫx��D�]tuM��(�܎4z�f���N����GoUw>�f�bND]�t-�y�M��;9���N
���.E=ʽ��}����R�P�}����Y�m:�ȁU�Zb�q�gg�c�8�`.�x��[0�,<��=�3�fb|�cg�o���v �`��is[�#f�D���ko�v*؂�-��uq1# �Jܷ6b��Ǵk�M���V�bؗ[�{~�X,K[��N�*�J�g��i����$�e�DOUA�Z�N%0�gFho�W�p�v�럐�r�n�S�]3R���wΘ;�"M���C���3�m�![yO�`Ҹkm���م0�;^��^�CkS[�8`o]���;�&_�o->�;d�N�bj�0N�3u�+�x�f2�{���w$��<n��,PsS-��چ�y&wf�v�l�G[����t�䒶�%X�ܻ�w
Ƞw��T�`Q<�O�g�@�ΩVf�D{��Oݕ�b{'��U'�,��������Ad�o:l�s�j�*�p�]xwI��s�w�܁5��y����`���Ht�㙾�;N�dLwP{�a�}Q8!��m@"���Gkغ���i��ֶ����*�d6������{Zw�gt3�ɜ
n�y��y8pl齨�0���P)Y��(���M���M�\Hk��Zy7��+�۸r�1�,�}9UG��Y��E�����3,�{S�jA&+2n�u��;���2+R1��TJ�(\*+��!F]�V����s�ϳP�:X�p�]1�b�-�ھ�2'	�U^Xr�T�n��s�x����^+�%A�����s��Ҝ����}
�
@1%�P��doj��3�:i��=i����᳧&d����r.a�5�`I"g*4\�kP�K|�܊��cup5nғ�Wqh(�Q�iJ���q�/nP13�S(��[]���u*0��q��e�5�U���]�����+��|���蒢g<.n�n���v^��D����{S�a���,X�Y4̗4��*�Y4��bFf��(쒲z�Hg��|i��}5�@FQH�j�㻭�'Y�u1U�O�X#S�[�X�i��v)Ήe̩�}\���UL��s*�_!���2n��k#*VuR$���]��T�o��:�3"5�!FD���}ݦ�RJ���w��R���D��Wd��T���`b�B��=
���]�X\����Ӫ���}�qT�N���8�F�q�z'с�G@=^�~�;�M�# �k+=s�s5�r��H	�Qkpfҥ]��n'|�(P\�jF<�;�Q0iu��"v�n��D�;0�p4u�+jsƞWs�*�h��F[jU�k����X(w`ِۚ��8j 7.2f�Xzo"gf�ޭơk�@
w��;Wا�WQx��wF�L\����rm]�0�nAUj{��upY��v�0��2��WgI���5�3�E�����f.�[�����Um����륞s6���'(��,EWX������=Z_H�ӛ��1N��Bv���u���}}M�]V��24EǷ1���>�bP�5Aָ����Gg�S�M�%,�,�f:�Ib�z2�r��}��u��O��v�GU����I[����O'J���$��)�\!YtN���k��h�	+����ê�!	����bnbr�sZU��®�]Un�U3�� 틫�������7��tr�03+6����ή�i�9�L�;��"¬�n�F:ˉ�+��aQ��J�b�U�9S�LY�T2��*�E��)tt����kU�2���He�oD�;=j�ȷy���wl���a��������ݬ+.��B,C�
Ogo��9��0���d�Ĭ��{c6Mf=�2���|�)��{����7�kkx���*^���Nczt_E5k��Y���tN�rS°ㅖ�P������ �J������5T������c����<��Ҫ8"���poFe�jŘ:�Y����[۪ptl��6h*z�0V��%���V|��Y2*	w�ka���W99����j��ǦnB��X�LfQ��{PȪp��2�E�oA�(t���l(m�v#.�����T�յjU��]=V�%>�S�ul�7w�:�z��J^����+�}R7c�M�oO�[wȊ��Y����v�>�5з�QSk`��UR��x���Xڔ9űwPo#���FV�)�oB� ��5Y$/3��dv�O��μx��V�ūT7J�&�A)s}$t'�"��C���cU=�К5��D�9���2�\���Tfa�<�k��K�]�j0D�8݉#1�1�[MUD�bsy�
�bM�z-Yl 6ԌÏd���归3�\k�tԽˣ�����/F��x��&sue.z9fWT�`y�;}2nf3@̐�:�9�뀠��ͮJ��/v�2�d�&[���.lE`'2\���F	^#��#9d�0I�JuUu�N��#_��k���wx�brUJv�Y��޸N&*�]z����+��R���{�"�vL��Y��E����l�;X��xF��-�_N4�#��1��3n9����ݥ`nU.����LGJ�M�&� ��Wl.�U�ЖV����d�H�1�q���hi�`�]�k����=�6j6���HKreA��U�"�uז�gv/�U������ɝgUn<�&��gv�n�)��̈+���V�B�<vح���q��3w@ˇ��꺐��c���Ro�w[�e�5�ܹ��
��b<����\/:�O������k��J�P���2[��y}�7���Ved�ե~޿`O:�8�����>���s9״.tS»L�їFw(M9]O��BP.zn�ⷵ��ô���]�����d�xLN_O��S���t�قЌ鍌��Q,I�1]F��Қ��ۨ��.F몫¶��_�Ԥgp]A�����L�3p�]��ʇ,]�[��u�Ț�ʄs����N�����%q��u�TD�b"3��7ZV�U��$;�ccl�b��jr;YN�\NV���9���6j�d�(�X�^����Tˎ�Z7M��t�:*�ݾҺ�����{�	k��X��w<Du�0�0���4�wNM��\�6�����Aؼ�����`3��w˘�|Ki23��4U��q+��4h��P�M����p{9$�v������i�ԁ�h�4��U����.���P2|��y�幗���ڋ����hX6�·��s}��؝g=;齢�s����ߝ��l���H���i��u
O7Q��c%@���v�C{隀��*���sTbo0Nu4���G��ɻ�٪�uMJ���fa�B��y� ��8��ܾ���S�hG�գ
�j�R�iכǅ��'�&��1��;�=����2e䩹�U/� T�����=*yD�uj�nQ�
�������E-��l+0��b����l(���'k�n� V$F�s>:�3#�C�٬[�Bk0�y-9�y�ܷ*�3��I�4N���;}s�2�dEi���̾�1*B��ӳ�,���{V�d���M�ƮDzgX��β��b�z:ru�s��p}���Y���2-�y���B���N2�܋J�d��e�c�ķ�gWo�t��JR&z�gM��s�u\m�kނ��p�0�H�U�f/O�����;/���z$]z֚�V3�T\�����"�c����m��S��|��O�nk���e���gcDm�2�ug�}�	TU���m%&�� �g8p7�\�7SyƋ7�(��]}��511����:��]�_$n�k'iԹ!S��AF�mþ�U�.�ky��V{�./�I�]T�u�N�'f�� ��Tu`���c����z�u�Ց�U;�xc)ܫZ��XJV싓Y�Ш�;1�{�D�hv��]�qD̥���j�,H~t B�t��y��[˱G<�2�cq3��3f�j����^m5q�wF�D���g]���PVn@�0��B�bn'��-���wW�٣e��M��e5���;b�]	ȹM�T�l�$�V��C��5P{�h�Ε��d�UKw��0׳���ɫ��.N) >����*R9�"V��>٧�
��&o.&E�qƑ�Qf7�:�8��ع�dj�̬����A[lNxE]���ӛ�G?(���䚝��U�<�d�{qk�Gn�QJz�.(6L\o. J��U�`V���E�\S樮za�:�j���&�*2��0,�|�&9��s�*5E�amF8���/�����P��3�{�b��W��8�Fi�7}��(]k�r���f�lr2'z�7F\k�e]��u\j6rŗW!Ը�p���P�8��K踺$T�lz�nt�D�J��HYo��Q;�C��Ɂ9�e��Ej�[*T�\;5�9
Q�9�����ղ��llg�2�{9e�����W}zxC��i�c*1u�v�t��=ӹwyX�eؗ�$��1����ɋ��X�	��R�F;9Ngeb'f���"�]�V��7����ȇ�q]����
s{����3w�-ܵ;ٰ!3�0�g�v=y����zB��I�l���O�::�����y�2�t�稪�w�W���>�uI�=��]���ˉU)؍s������.��&��-ۻtt����vup��1@�4t�О��F� �
�&�S4&j3�q;n�)ELɎͭ��UѰ-W>�5�\u�M�s�mEq��<%�[!ݼ�/pؙ��ۚ���u�z��\L�oD�6�v�%p�)W����n��ȫ�R���5h�1��-�O�J22������%�ٌղ�]���U��U�!��jE��}�TQc�6] �C22���dP��GeK̻|#�2��#��0��ԅ�Q53g����cgaL.�0���M8;(,B��7ky�n��eǔ$�id���k�T*LN��;An$�֔i�F���:������|Bɴ�R�ZA����to9�-������-	}S�ٓ΢�]���8^I�b9��+n�����``����͞ڝ�[:��X]Ժ��u��if�b�8kU\����qj�F�LJ�qK]�S��0�Y��������:خ�k��ٛTSk#�R���?Mx`;�;bB׵R�r�b�Ʈ�37�tү7k�fゥ�r���O��]ǭZ�����sn��k�o\uc�֯cT��4\u���{��| �4�+
�LM�.���kR8f��}��cw��sԲ�A���ޣ����5�Odvl$�xg�,����G���k�-u��+��'&�̊�w26a���*21c�|wL�,���"���ob$)E�55���압��ۺ�DM;\MJ�m>�0i lvN�|�s�	�SP;u��ށ�s��b�T�*x]յ~�9ԣ����I��ʍ6�7W+܇��PI�Us��y��]8.�]�֢P���tN�2�F���OT>����Q=�yoz�C�r����[���.Fku�c�{�u����R$D�q�3qf*i��}�ú{��i]����|;b�x��7<3�֓X�Ed���:�#�uM�5U�	g�� �NP�'Wd�5Fc���U]�n�r U�̻̎�sKjVH;ϥy�s�:�hU����Df�P����i��ė��O��l(��@������]�f��1�mc�R���ei�=�D��%{�l&	�HV{3�vrl'*�3q�z��a�@�[f���{qSKKfA�%��~l��P�;U��\(�p��r���.��}�5�Dzv��c{$Luk�ɭ�.ܧ.R��7� ǣ�7��F�K��m�P���
2�Y�˽�`�)�=�\����I��r���z�1i��霮Q!�7`�;��j��������kA���wg��D�5���x1����&Y"������t��=�
��i�s�ͥ���#�	һ��=�A©c�z$f��������Yw�2�P��2e�]�v6h��Nd_JK�yL�/.�\P�eN����\�*'��u1s��zճh�#��5�Wq��yͅ�Rh��p꼃@Z3�.�g�/}�SQ�(�yQV:z�кR�Y�h�NE+&T�\hu��7e6�k���]v�.����/Jm��t|Q�Җq�%�Ý0�U{��[��*�w�v�15}���B�m3X�U����6��SrG̛�}��*ƞѝ|N�9K_\,�bc��H���0:��9��]Evvl+�$H��s�U����ԯ��J���D�t��pЕ�����-�k�Yɰ��aU��h�9���h�ҫ�#V�:C��uV�8�D�̛����{��Xκ��^���}���S���T�[*�w��&:Ҋ0�̲7z��Yg��/�J��9V��E��'�ci_�+��V6I��Y��wv@�ۻ��N>�.��n`���z@��--�bj�W
r�T�T�`4�"K��{��qu!��Y.�6��1]����1� ���:Ӽۉ8W��.��ۓrqqu�(��ث�8�u;�P��A���k�����^V��}Y�#uǠ	p6�H�dl�ڊ��6�d(���y6�u��ˌԪ��fE�4]UED�S2�MN�d��,��CB��t�n��1��f�wVٔ8�w�5TI���c���:�j���Я6c!�M�lv�	���/cU����Iާ�7����v��r�z��4����͈[�P����nT���sr�oE_u�g:��'s�jN��f��dr��Wq�s�چTK���]N��\�y��ɚ۩��婶�d�s�͘�oU���	g��	�,w'�*�t���i�~%�*�7l��V�{(��\�r{�z�3s�+�t�[��Ol�����F_o������tS\#v4]e�������n���8���M��82��:ܢ�&��;k��S��,��o7��t��9�`���jf��Ԧ�.�(-��}{��aҽ�m��xCN^y��Nc�9ʳ$���;Ѵ����;�f��6n]�Θ��i�LM�L� ^ő]�^p�ݬ�T�:�N}MR.�k5&�"������[��b��eY|�=��lf��X��;�I�V�\�F>v���v�,�1𩲶� ����{
�x�hnKN�u���2�z��

H�+�zwdˢL��m)�"����в�7Q�:��V\��������i�ccaVY7I��;�*׌���Tj�Όw��*�&�M]��}}vyke ˝��ǲԌM`��Xf�(^�x��Քd�jƣu،�N����\b�U�=XX�7��t6�L`R�����([�'�v	�/J�({0�=�G��pI[3D�����U������6���#�K%���M������צ-�E������Fz��ť��>��i*��ϯgj8D��!��g�	!�����D��ᜦ������:�H��d8cFY}�8i�eʌ�_��Eq����ٵ5s��GU{����5i�Mڤ6�s�@�J��pMP�)�s1[ uY�\i캍�<���`݉�B[����f�o1Nz8edt4�����s��d����z{vb��٘�]�ڊ���ٮ��9Nݛ˺Ύ��Q�,�9�t��^������m_�9�}T`�j�3�[�6VuT�+�ٖ�jܲ&�v�wnٻW�	�Ge	qk�����Gf���\�/i��3/��6�D��ݵ�;��������UE��-�����ƒ�aXC����zg��\���Ƈ�w^D��R�y���H��n���c��呼�^����b/�*�l�@5#+�aѵ�>�pg���6�6t��$�U�n��C-���c�'�D��=Z�q�4-Z��#'v��0T�c����$�h�12/�k�� �S�{�1�n�\�ф7o��bۍO,W�����@��=�8fJ�"��7�3��qlœ=�ܞ3��gD����1�;(�fˬ�1ו���a�UO��]��5��z��|a�r�.��ou��4�z��2�񛽸�:��iOH���\wd���:������%�̋���w&�6�x.�S�Ρ"�M���pu�ݜ��;lUәO��;nk:�B����e@��b8�IP'��i�0�]dVN-����w���B�0X�-����qŔ�:z6�`ݓ14�Dv"�/���2����Y*��r����m��ڑ�Cr2}��~]��{�kY{bǱwO	�4:�.�s��[1�>ȫ�|�z�]f����z�۳D�2LuWS�K4Ud���"�g60h3�f��5��r^�r���&�Gtj��x�;q,�9�5'v�P0�ٕt7rQ����L]�N)����$���x�����B�q1w+�}C1<ѝkI��NOw��{0@0�)�\��>�o�C��Wڲ��6.�s��(���:�^������ᙻ���]Zk&�����3��$��3J��Ӻb�=tV3o9u�n�p����Q��h�BݚQ����	R[S�a�iF�$LH��+�C���,��ê_m�o��*O7u�b������f�;��u=�!���j�mE�t&OHx՛3#Kjsn2eUU=���MX�}����z�Ѯ���X#3r�*;�7"FɾȘ�{�ʧ�w��j���TM�wk��ã�/:Nf�r��vvT����<���G'����cEm*���9iLP�R=�%.|����Q���8ʃs��7�Nu�ѷ6��j��]Z��U���Td�� ia��3���u�����.k]ٛT�)L�����E>8	�G�Fm�<N�A@LN����v���MX��uQ;]�:j�yY�tXW����㦬	�ǚ���ʕ3}�?#���-��ɱj褩UJj���fڷr�˙ݵ�M�W5ʹF���sI�r��ncJ���"�k�+���2	)c�[�W5,F�Ӛ���r]�%��9.U�\�lX��W6"#c\���ŉ��v�Int�����r�h�ݱ�aVa��A�9�������5�� ���~���?�=��g�c�j˜��I;�T�7�'��?d�
6�W�}K>_��>_�b^�#���m��Lcv�N}��~:��O����/���(�
+�`'��'�;e-�?-����GB`���:EP���Ͱ��;��>�} ���04C �C/��;����
��'�7%�ˉ��!���ߎw|0�����%�����$���g������7���J����G{Sy�g�3�=J2��� ��%��"f��	��b�����#�iQ���t�w�Ԇ/�KW��*�.��F�����3�V�S���
�nє���^��Ƣb�i������zPg��-���aU����Ciz~ƭ�?9���Ҟd/U.[ �wW8�f����k�_3 �/�;F�7%dU�n�x4Uf��Y��N�Z���M��gˑ�L��/�DΗ��|����	Ԝ#���:�J��LF�R��#�SI���ݥ)zl�I�vAr��G�oC�ֱ��p�ͅ%���»�ճ��^��e�h������]�W�?WWa���a�XQ�}˜#x���2��lRR�߹�$�^-�\O�-��|�b�ѩ�'�??��䊯7<�2�/2���g����5ax�-�Q��b馕�������Y�@v���'��G�W��C{4�]z���pA1��;��Ko�����Ҵ|�y��ݵ,���9޹�*�EE˹�ДK�Q�V��t�%���oN�N�!� "pV�����]^�&Z��~U�시�{�غ�l�Z�g!��`��`�KԲ��۝?��^�qfg���9�A��f���F� �I����*�����=*�p��.�R8��<E�����20�8�霱]�ev�-C��v�;Q��3�l�OV��]3Ex-��w���������\{��-ZT��Xx���	��Q���2%�'��R�%��C �xV��S�Do@��F���d���<8d�F��'��g�xE�7H�A��dNj��i~[/��\���{�+�����8'�푾��Lv�vW\�?��Zv����(����k���Es�t(r�s��i	�S C7���X��c���N���������N�a�^leXGc�P�"�|�d�[���\�9%�4)�yF1Ir���2B�f�dFi�K�g�w����*���\����$x@�}�#��=l5m����8�F�7.���{L�P�dz�>0�5�
����}�j�I��9�#e�ɩW��V��ZE�k-O=e����tW<Y�o���?���m�4s1�p�����j�X^$_s_���W�{�r�ur���/�	"���n䮣�ܹ�_3⧉<R6}4���z/X��_pL��J�D�4ި���<�Sψ��B�y�x��-qt�CM��[|>�Tm!�jO�ĭ��A�NW����u��ْ."	�F��4|��6�=���x^Mvt	�ZiH�b�)�kz[�������(�|>�>�ROd���_n^ǵ���{PLU�{�������2yVV����H0��c|��.����Dv~M��B����(��e�*�O*vZ~���?�&E��'���޲u�V;B�p���8{��q)n�b_�����9��x�̔X��Q!.̬:{�y�|Z���w��k�@�ִ�Ll���@�G�Ii���y�y�L���(��]�Ұ���t�wx���4'�
�~ƨ/r�L���V6�R<�Z&mުC��CD�n$���-y��d�@*��=~��&Xؽݯ��k�S���o�ӗ׈���^N'Lj�_O�_�rBL&&{���k���
��"��*��\Q�v��M�Ҹ~�!߹+Ϝt̕�oH���fO����0�,Q((���:G�+R��b��2R�Ѯ����3���,J����c�}��fW1�73 {�T��;��Z��<��1@��T]�
�B�5��E%��z"�;3	9.��کE'XQ���/�R�+�g�A9�W8��S�|�2S�(t۲&���C�,q�$g��r�{�T�t1���]]ɲY���j��.;�~KL=��(��5¼�����y��U�\���j�Q��<$�u7��lV/��?'���>>g���/�� B~_Go�h��S���6���������w��?�֢j\�����S�Wo�P��_���>Q������n���klOI�x��C6�ߊ����ܴb�+&ݖz�@B��~�o�u��xV��������ϋL��f���!מzם����-�ީ�iu����;kw��|q�-�a������g�f�ݘ�Ϧ�ݼa�q���;��Lg]��4oE;��M��F�Wz�P�	/��զqW�\�d�KJݻ����w������L�Hj^|�����V9��S;�~�O�tQ4mAz�w���߮Cg9������i!<�V2�V��@j�]���o�y����J���o^cYӡ>�Un�+a>�������k���y�]�p_P��ǃ�'�jѴ��������[�/�R�X��\��C�*b��^�|x�6�W�`o�6�MJ9��I"ʃ�j��x�.�N#�^��W�mύ���`�g8 p �+���7G�"d�����y?��;��=�Pe�>V{7��մom�q�����|س6��(A�@?���>>8���B}�������u�޾W����߸���O���L$���{��>s����W�a��bg�m.����G��+�����[�\"g�!_o�H�r���9�*��5w�<Klz�;�;d�"��������fk�N	PC���"F~y&k�o�O�"8ATWrר���A�1;͎!C�[�k|8}q?�:l狧oP�	��ξ��"rN�̅�Ūy�C1�n���!��WuES$'5�����u�=tx&?P��4b����f�\p��&����s������ac7��T�����3���'k��J�x�[���6b{��&�O
�t�C=/O�WB$_���P6qRb��v�1y��}2s;� �19P�#G��UL��ƭNM���n�#��?�ă�:c�Ҵ���LY�n�^��������EwfI�>5�dVU^m���LZ"��vXb�S�A����"�_�B�F�޼k�!���'�J$�q*�*MGm3ÌԎ=-J��Z�m��b�5Ȱ�WRƶ[)q��8�#����B��;�w�U��,ۇG�=�IB�E��v.
ΐua���Gc������P;V���2Q��I��>ދ�S=W���^ ���K����(��.4�t��.�"Q��0嚅܊*h��rA�@�̸B�j]�����[��4��B��.���K�Kh>��Ĝ8����
����6С���z�D2f7�ᐭ��M!5,�Cd,͢ޚۺ��x`8�h�Lw����$s.��\R��,	%�Y��#��ƪ�B�+�D/�����gd1�uVIPg5���Ю�y���.�z���?����	�,t$�����6�����G�����Ţ�0�Hcɓ~�cӎ�})�7� ���0��̤�Z����w�E����ފ� �(dI��°o*q\U�ԛ����v؇Ԕ3y��Rv%�{.@
|�:Z���.���o#mz�v��Q�y�h+9���^�sH$pbi�]����9GWc�#����o��6<l�gzQ�yq��m�5�Z:�]��d���άL���&TjW_���O�nV��y�Nǥ�.ZՂ�R�%��3[�����Ú�I�����C��N6�X䐧Nї�6(�Ȇ<�]�8����%�����Q��c;X#����W0��r��|���a�^⹮�R?h�?Ũ��iĔ��m/���d"`d���?�e�D�p�T�����M
Dr���!p���\��c`�a9#�a;�=����(�W��i M�������ַo�95�3����K��K6���)�>ݏ�=��c��yz���T\�[�[���ށ�=ӻ�������v����̶/�z̈́d��VSK,�K���d�e�ԇ�L���U TQ�%N��*�W���{DkH�������t!�erN�nQ���쨻�W^��� g�R�D�H{�� �<.S|�������Өk �w2P���f���8�<�F-4��S�M�0�TjQ�o>�����k�I�K�db�n�kBue�I�5mx��{�峕;2TR��&զЙ�'̶&@�:9�Ҷ��l_�go��d�h|D\h�(�����^*m��e��������j�Q�no�(��јQM���8��F�U	1LX���u���W���ˢdF�́��#!j��<�����#ӯN�[D�j��u���4��!{-���WRR���C�����ɡѥ������$��u��(&�Dx��-�Px�1�2w��r��*VP���nG��Q[�Q��2@	�h@J��]o��4rN�x��Ka Kb1���"ҭ�_�+�eľAf���v���dj+zT��}���\�"V���y�2�e�$Ix�W��Z�B!�ps���/���S=|�l��&���?n�"!�NӼ��0�D�G��3w�ـ������"�^[�qt.Bn�g�,6T�ѡ.mB;n7�	7�ԥ-ӺV39".�]�[�8��?EK!� �;�s#��l80k*dsǄ6��-m,��h[�mps���������������?ݿ�~�+4�/�_1O�-ݍ�7+����c�F��U���&��m�~���W���?�ɟAT��:wa�奮�P�^i�Z��$�1:g!����+�1�W��g��+ry�ņn�|�&z�!^[�i��袩�oߌ�D_������ۈ�ş̴���V4�][�L�6���8�/[�,&�r�=�ۮ�����X�X����Y����㎈�x�D��]��7q�����=���*�W�xY$y��������ؗÉ�A)��/��];�n%�H�ԇG�:�#�;��Y��M��c�F�{suը����"���<G�>�IF^13ɔ��ӎ��Ή<�{v�T�51����C�"^���V�������Ü�	�`D�1;������~w!�^{�>[���7}�����z��j1h����<��{����K���j��)� �$A. �v�E�������! ���,�w��2�#$�\7��G��ȍ���8y@�~�Gh�8�E��3D�l�Zi�Vz"�Q�k}�X�˴D�zMC �����~.v\H�}��-�54��*oXo�w�#-���o~��ou/�w��U��y�x���Υ����Dᘂ..�����j�q<�!x��3dkd>�|]���<��o��{$6��v���JQ-Z����Fe��)��(�������� ������O|�Yt(��%�}��I@��JQ��o�$l�Z�YD@+E���eQ����a!�'�?t���Nz�2,�}�X%�t�������?�<EN�r@W�1S����������E�"xZA0T�ƺMͶ���K^o���2�<6�ѭ�|޸fZ���ǐ��!H�!B�HR! @��9�.pp�����?�?r����L�����4��'d��⏼�oh�)�J؅s��$�(�!0�b�_z��P��pa��0�,a^�I�|b�s��8`֢��"��Ex�=�� ��5gf�iI��+�{-Z��'�Y$M�T�J�W�ȡp�R�J��-xFC�,K�Z���P����DR�g�q��$�lR� ��"��UE��	��%	�Z�XR�X:��'[�F�Ԉ�P�oP���HMq)���1<80p ��Ȥ�`=��}�����y"<�C�� 8xq�������ʓ�UX"��H($�X�`�# �\������7�{�(O*/��B13�&�T>�����PV�ptu�B�N��D�n�48�ݞ�WtӘ��蹞pv[-��h�ܹ�I��6�/� D=��s#(򹻡Z�Ǜ ټ`i�$�����"IS%�luC�`_ruy�]r������� �F��g�iQ��q����8 �!��y��h��l˿����t�f�d>�ǽ<_f7-�n�ڸ*�P����mw���}Yp��,}�x�﹉4�O�/������=/�<�ς{�]�_OM＿m�~��V�޿=�\}N�=���I������n��֮/�Nʠ�{����w�6}f��WDV���81}��_��?�Y�����U��B'��0�O�p'*D���:��bEQ?�V4q1?Ƌ$z��Dw���~퇺�R�$Ä�)p�ʯm̠��d���X""j�
E�u�|HmBcψCO������ �T��Ι@����ۄL9�ع1A߫�w('���b�ދ[�	���r��Lsl"�A�L�\i�����G�d��p~���a��A3E-~��`�w����<8Ҏ��-O�T�G�\�T�mu�r/����*��/�����@ܰ�Z��7�PP��g�&mT`ƨ�Eٍmd���U��J�BN��A$�؟o��~k��;R)����o[7OA�K�Td{sM����pB]�!2t�{�I~u�T(]:�4m�8V�'S��l�r�*:�:���%"c�T�&B��#�/��[�@�n�߼֠���H��-ww.C��xA=���}#�2r"%k�ьb��xD=�t�*��Iި�k�;�-�����WP����Q�!ήp�m�wft��. ��� \�F�-1�(����`C ��ɱ��ƆSXE�N���6H�9�/LX�3�0q�'�ގ�M��>���G���"D� ���K/%N{����Ž�A%��N�H�*��#+����w\:�1����I#�.C0@�V*�B5��I8�{��0����@���]rM=�^M���'�0fB㝒ĒA��s�F!��:���ʠi!�"ɫ�X�@��/��gF�`�B"�1��/�͒07M�n.�Q�Z���)a�:ʯ�V)�����.{�Y���:���E^�E����EB#��
��~ŷ��*Oُ!.hp]���z���.;k�>�q,E� G�Ƥl��ڈ8�G��s��S�^� W�aqA��7K1f�"�*G����h����i=ےAu�j�|$	.c ��q�!{Đ��/��+"��7��"
�R:InԿ% 7J�g���Gl�U�.0TW�F���*}��F�%����'��c�C'��̽�V�0@Ȏy����yb�/A2�)�o˼�X�U���S��==���x7!a�����d�2�B"�*cr�J���7 ~X#�Fﰭ��V��T:%�*K�qUk�ͦ���Re�ikW
rSõ��ʑ�]��]4GaN�?r��/�<>���*쀲�_>v�xy�uo=�{��H�����L��5*�C���7�z2�J��eDyp� _\���b٭W,��	
�$T���o�ĉC��{R�t�I��E���@�^m�ډ>�T�M��"L�&���\�����ej�T��7�u�N#<��/!�wd�����w�1�dP@BA��?w��2
��W�\�I�0�t��D"Gi��i��t��+�%Zs���>�!o^���8d�G��_�c?k���5��,�I�E߳��e���l�����Qn�\4�!�V'�[��:�}%��93M�HPA�֢�H�C�Pb	������Z�����R�n,
��F�(8�YQ���):�-����t�ytz�g�����~��: �����ܲJIQ7Fb����U�"�*$aVE���A�O�:��쑴?R�6C ePU�z��P~���4��5@�������Iy��W�@)	Z���\�T��'��c�0��^���살@��jԨ����Shs���hH�Yֶ�C[��Ya%�:���>s|�"���_u�FpgL^�H{�m�Yt�t�C3���L�7��{ OHw�=����x0�3��������Q|�����������`������#�{�������.�u�̈��T_E�aN�>�ϺnG��J����4�H�H�Z](����f�����,�j��!+��s������v�T��(X+ޢ�-?L�n*d���\���wz D-�c��=�W�˛��.�UU0�4�	���>E1;~�Ϥ��	?��3���w�]h�Ѕ�+��/�f�>8�(�O��|�4��	��z3�Q�G�oI�b�2d��_'���2�!*�����5��뀐��������jP�"�̉�b�v�?Q��AGA�[�}��C�^l���o�)���;"�Q����'�L|s�Z;�߰G��n9�~�[er��s���"��(`֕0������;��tB�����薙�$H;��s�

c�ܭ�5n���r˖�t����h�q�f�Bx}�Jޛ0}��Y#E����Kg���C}�f;V)=ıF%
ױb �����=m�x~������m4���2��SJ�5�X�]f�0��M�o�}��13[<<L(-��I���X#�z0�9�i)'6�E����_J��4��p�i�̒$a/��� ��E����63)e�]��mu2��A(>߳�=I��Kqm��BH�w���L����u��.�lf��m'�(��F�����k�����ƪ��q��I/3�^��1Cz�<���r�ׄ�`�R>���F���#�(�Ҳ}=Nz�ƌ�>�����DcDD-0M{#F*_p_�O�̾�0�:ϧ����%�츂�I�����e�	��%�eR'
���;E!���N��K�cO"9��~���#�^�W��|��c�M�4ڸ�6z��Z�̅:=c#�:���I#�u�KHBe��u��v�k�&՘y����(Y>��~l���0?r
p�߄�5�J�rx�Cr��,����B�P�c�u=E��Q��+����t���kM��ǯ5�~{nϴ6TG١ �Մ;4Ğ$� �+�p�K͞�Df�U�To��C"NqI�9n�]-�-���0-��;���$`y�j���!G�^�c�h�hNp�(�����[�[g;%Zo�2jv̢
h�2xҰ��_��W^�H�O�U��A	���ЙF}j�ʖe��堧�[��mz^��=���=P����!�~9̧����T=��]�`C��%�eݏ��C��X�&e��9�z�S����oo�Y2rz�s՗(�Z~��\���9�^�NF(��`�����Kĸ�K�x��2��(bԊ��1R�x�kk�Ocg�$�*�L�>QYL,^���i`x�L�6��Ѹ�[�;ʭ�E�0K���KٳG��ߤ3�p�њ�2���p�?4Q��ͯ{bx{���������3q� �0��"rr��6K�� ���5�[J9&{���@��1�3�[������Ǔ�_�_hĿR�H�:������9E�"�H�{B"��{CP��YU�h�&���]\��XA�s������g0	�W�mG�6J�Y���B��C�*�E����B���jkd���[�RV�d�[uW�@a(*���j����ݖ��~�l/�?b�=�}�l!����4i�[u��t�,��U�ײ�1|ʘ�p���0_M*���CUa[bas'쇜bEb���˳���1�����z��ϝs�RzZ�6ɭ?(木���GG����@נo�?tH�D��ߘ�&*US�xm.����g��~d�6y3O��x>}|�)���8��4�H"[<!L7+�>G2��]��}\G}�R�e&�"�U���X��6�r^��mv��r�'�x������o�;�]ld���	��5�I�G�C�gs$�=������qU8��D얉�]��h�T�z�S���Q��YM�`�ܦ<���W�eK������8�]�L`K�.¤i+d�:��'�����ʩJ��HCN-}���g��~�k���k�X�mO�,� ��h@l0���V��gj<&�kF �4eD|k��ǫ��=a��UM���MT1��c��՞	H��3Iw8���A��(��þ���7�d���IXp��Wh��n�=��ݫ��|���ca��g�I�'��q;d_���.+��MBbX��&���/bmqz
F���451��y�^�ej�i�)y�I��z��Ш�5�8��;9���F�2�D�A��X�οkg�ħ��rq�àu`QB}����1����)r{B4�D{�2��oMߺ|�@K#l�q �j�H#� xM�2ļ&�|�����<�������d0��b6og����S^�?��j�r/�1���X ķ�
C}/�mx��{�'�GmF�=n��i��5��$����5��n�vv�/#�N�Q	��c��R{����?T���QL�)��=U�J@�T>��V��~�ևUj�Ab�A
��#U3T���3�K�FU�?��Y����G�!\�n��;tp1���֨�������o1j��E��@�M�F$M���@�6��(����EX*�o}6�#��R�TY������3�c_^k��seL\r��åV2
'���%���v�Xl�g��@��m�ݞR �3(��lMy�w~�D��z�
<��ଓ<_-Q4)1!)����/J~vm�X��JA�B�����%��v�|}M���\~��>O �q�Ћ��=��JQ�;"�²�"��G�x�dM���Ȉ]�`҂q�7`���{q�#�+.�x��ߗ�Y�w!B?¥��(g�wC�Db���JW�y�|`����W�:c�d���9�th��x��~��jʞ$���(��m/g��|�̳�(핓ݒ2d)��6��{�۴�J��IGr�1��u��K��x���m�ggm�� ')�C1\z�-\b�I"�p��*�==�2�v�͇k��~rJ�b3���{���k�����$`n�2�@%{_�:��7����bB���M3�x����z*<��0�GjZny?���$VK|�Em�jwbS�n9~1i �"2Na���;��d����n�K���w�n��)Ȇ�)];���z�Q'ƞęm^�.µ�D�t�~s�KF�om��N���:XdM	A�5��\�<�(�Y=\���p�4[Q�)�����b��G!Qc�Xn�a�=?� � ��/�<�����8��N��KyQ���Q�^MX�/nҲm���\=��-�(f�ȇ�|EP&b��{x�3D(T��Ù�R�x����[k��z|�$b1'��z�6~�(�W�l�/�^�J��;�x��#b�k��apF� �
R��.�z.#[lxh7n#c��%�"�Ʃ��l��i�P|6�����d��|��55��|?��� �����7^��#]�� -P�Z,ޅ�M�<M{�Ǽ{�/gھ�����s)�N�M�>Ӂ�WLV�&��"��o�Bށ�՝��%����v�["]�\`o?i�w".�U�&��b��l��"!d]-��=���i;�\1
I�H2������U�9�8��SY)ћ����5��>yõ$��yZ�r\�z��L�	ڒ�şLB�J�"���XE�+���ήEueƥ��� Ì�D�Yv�i���p�o�:�:��-�A5Դ�2/G���A�2�l��0o�Y	:'Uv��GO?(�4�ݰn���Q�D$��_&�#"�t��(���H@E���矉$���L�D
YE������+.��y�ÏO��ݻ���<&�*4f�u�?��	(�}�$uU-��S���9Ӌ��Z\�!�UB���1�[�2�7��s��<d,�!(>}����j��|�|�#fvqe@��ۄx��>�>���m����@b��Yg��fք~Wcб'dM����/�
'�	x��/a�Q��'�$��i�����hR;���&����Ȉ�?,����侈��nl=o����^'{C]��9���k4�
i0YY+y��D`�v<gO ��i�b�X�0vi�:"�^����Y͌�2r�u���DR�̠ J	����n��!���m�7�)����",6lKWY)3���M��d(Z8�D)�|�o=>I>�U�ʠ+L_���D����D���%�Χ������"�K��X}��q��X�e��ږ�܎�g���	�q�\���3�8�iv��dU��Q�))'-j Ѐ���ɘa�?E��Ϲ,R����=k�t\���Jr�<uM�v~��!C�h���U�Xt8���]��<����F����-6�hH�;��p�!G�d�y7cY)��em��32,S(��/�&�_sp�-k�yw�?Y��]��k
;��%��eH�z�Љ\^
K�5�k�|�R�P*8!�uy�B��!��O�-���(��S#{�3:(����(1z=Y8�)��1ۼ</���_]�rs�i��w�9�f���ߕ�H���P3!¤Y*�ך����$���˴#c��݄	V���
��]��x�A<J�N�̞Dca��I3���I�R7Q�LO���uk��gr��+��2=��NT\R=�ˉi�C/��~��13�?�.3ի�%� ��؇��Ns�˺��1��pE:R�Z�$��)�����Un���9B\Lt��U(�C	���Sײ�^�'o���bOdA���[@v�*�.�g��BP�New��w����D_ΗH*2��.���>o}��1���s�6��h#��$����bT���H��>s�>T`�C�{Z��GG��ݶ����������7��2��!`S�f����x��8V[�(�s���)z�=з>��'��:}�sxW�#�K���ˍ����ތ(�8������h��$(0n�	|�Jh��Z�Ora�hJ��e����J!<*L<�Z~}�֒��x��Tv�&�ly���j�>ʈ���ۘ�l����Ga�c�%��g������=?��<�È���v��?M�ϛH�����&#�����Gj�N�U��-(V /kK��)����l�!�3�h�b��~0-l)r�U�g�?~/�c�����vo�R�@��=69�T� �]�����>;��B�#�.\h��v	�λ���p%w���{���+��ai�����bv���_���&�se3�BR}�G��翵D뎦*	�*,����۷��)tf���Z���P��af�t"ɒs�O����kf�|�oz:������M��T��Rw�8_x_'dvP����<�4\���_*4B����>j9��eP�B\Q	Mꔧ���7��K7�L��Iǫext�ѕ҅B䤨p7���*�A0C�$����#�r)@Qg�*Zj <��8�o1��?v�(RH�*#��yQM?>��5w*%��=zP���7S�(
�����"AE�
9{ǜ���ޓq+;f\b��_�1��E
^�h�E[��U���Q8�W�TbuP�&|*L�.�m���%�l��(��t���?s��7�V��7t�[\��5���9����B�5��r:\	�OP��OE�3׹�)�L�*I ��eIox=��ݦw���
!�ߚX�L��,�ͷMw.�-�C;��l�����|D�	��� ��L+�I�o:^�����&��pmTr��r5�z��T��:A��	V���E�E���Bi7�e%�@Q
$Q��{o&��@��%�r<�]�C¨U��|$������l8)wH�T�@�~�i��>��N���J�:�:�ز\?�I0H�ެ�RhQ���s[�"sC�w.�$���:�9g��mr	27����㼄K��`��ˌ�s�ۚvz��_�[/^�"Uj"L�U��5������* �"�e}h'}��%<�0ElI5+vDa���C�z���H���(������n1hG�_�)9іy�i>dqx����:���u����C+��eE��.R�/m+9�⴮���V;!�X���og�8����m^$2�ķ#DT�U��SaA=�Jm�
=���i�@t�oEAY��?�r�U%Ar\�\�l��(r�D6FLk}�63�	��k=x{�P�da�5��,��Am;@�>���,A�S�|�)�?���$��f���TqGu�����5�*>'uu��Z�BY�z���Ǯ���}xF$�m*���5��k]����^����n�.p��RLO2��.�������n.HDOZo�B��)� �$��tu��J��%>�&:�?�y.�9`�!!�g�g����m���p�����I~��+H�<ye��6�
�ڨ�ʄ����h*�G]�f{6�m���G�8]�_6W�B����se_Io5GZd�B������n�>��Z�dQP��`�W����z�/��!)lQmpw@�D�h)3z�>�W���
/ͰȈ��¼�3��&�9A��@�q5<���[Q8.r�xuK�"ǫ�ӳ��Y8�WM�z۫�Y �m�x�vQ�L�!"";8����W�gn����?]"���K��=������x0����\^O@�D�2�I	�Ann�� \�TA������O�2~j�;*Q����)�'Q��M��91"'���`��K�J�ϊ�M�����ڴ�$A	��������)�����O-�g<�((K�X�_ʎb��A��A���UJM��'�YO��Z�IK��+�"343��$�ety|���g��Q�� �T_:c�,��JEu,�M�;��Y��;�W�hp;��>��	�mK����D�`��i*�6@�Lz`�7N^��)JD������}����yz`�<�kr��%����Й�Rx
�Q�vs.��
����G�ʅ.bűj��bʙ5t_/���a*t���P�J�T`		�f�E��*��u��>BV;� cC?����>R�«�ė�<��`c�� ��w�ܳ%������DOޛ�H�%)���������VI&�m���7D���+�л
:l�\�2�<�Y܋~�x2 �J���ýpϣ���Ir�.�o��,� ��&��%�Z�E}wX��Z�ʬ*b��m{{E��~*�o
��D�^X��+�����vGZho��� �sOޢ�~�����M���PE��r�C�7�w���ھ��R�!����f��S�\�"NJ
"M2�گ"����ϭ�4�Ủm�̅T��mk'�؄3QUB�Y������A�p$�3R��R�ZfI7���9J��!�4���m!yx��k���3f\y�H$xd�g^�#c���j��Xpc�+0��Fe�r;��d�Ģ��叠����aC� B������G$?+ �ݹD�}j#eA��e���^vտr_�����}���0y��sO��~��('b������z�'��C�d)ؔ��R�� I.�	���;R��1$��D+01t(��$�챇x�"�6�`���!���z��%�>Ҥ����Tn�����-�[)�\��9��1�78���Ў1XF&�v�Ȭ�*LwF
dS�b�0D=��>����v�������Q��ڍr��C�"ڃ���;�����Gb���q�'g�P�DVh���c9̰SC '�ʡ�P	�R��0�U�X<E�����
E!�<	+���+|�^ n?�~�/�k���^^/����ߜ�D{�Lۻ)qj��J8��4�Y�or5!a9+�Q��HwD��()�Ag�/�v���WF}aɂ#�@�uKˌ������Hw�7��ܡֹh�iQ��"�v?�E�i��B
���N����{߅��E�� 4�H/h����6�n���jɀ����/>H���v��L(g���DD��ڏ	I��G���5��(������C8��ڇ7��3�.*7G���S�����IXz�GD��.EQ�36�

��۝�"Lv��!��{ڀE棣���"���������=�B��;�-*VF�@~��-�w��m�SbTI���W���Bޯ;q�ZVd��N𕤄�@����D��e��2�T2>��Pft�,���fLYk	>�m4|��	N=�<��N�(�ܲ��=������<����TxK�2��(3�m�̜�������z��j̋��aW�+��W�4zY���D����:�cG.mw�B�g�-@�q]堾w[H�6������֤���t�W�w)]�����Z���	
,:�� ��I}u1����[��t���W�`˶���a�JY�ҧ�t�uhO�F��yH�)�܄V2G������R��:ژ>�)�3��b�0I�׷o}�:q�od���F��
����]��i���;�m��4a�tT�պ���v��BZ���c4$�z�a��|[�S�W��b�g�U���
L��0���rI�B4ĳ��Οe��a-��:(��_�Kw�k��!Y�V�Z�s�g�����������z9#��m�|X�������K�'!)�]��H��ӫU��ڊ�f��?��)l�z�j^��'pe�^D��@��wOC^���l0v��+�o�R���d�]���7�T�W��2�\z�����(4�^R���:%�_�,���X@�Ҡ�c,��fB1N�7
}[�io����"�Y6ݠe�@�^q�J\�G�#g���L*�"*���7�3�tc/ӊpβ�����4���Ig[}�9yϠ^�����v�[q���6�!��VI�)�!�v�� ���w�;Cwﲠh�$7��P�O�>����(fA��,�M�J6H�U���w;m��7D��/Wj4f�a�͏&��eE7,��|�bK>%�iC��7;0� ����_�Z}�i�f-Z-��D��s�RǴ�9�!�{U��7��G��_q�7Ѩ�n*����7��JRڮ�i�q|��ͣ$F׺ʢw�=�!V�Eor��x�+����[Z�4vk�PMY*42��[o2H�m'h)�)ؿU5h]\�����s��1��,I"5��<-T�m-F9\q�c���%�iQ6��$#�.XuTd�1*S����ip:X��,|21�	����E""�z�"�%�~�_��a�2ѺX����JbO��RV��Ap���Y�"��q�6��#����.j�{������Y�X��iV����.��9��$�q��:d�N�6IEa�+�s��뽶��nEp�`���W�H����_s'��o�wA�q��M�ߙ�.u����ὴnl���X��|�髷y��8{r�x��&��F��պA�� �i�����
�$�|�(N�01Hl�
� �q�'Aͣ�.�C�E������^m������w�gJ���z��o�x���i탨.T=��9�+����-�׉kdڵr�&P���j�G���%�8���)N�Ӵ�$9��Ibóѕ�~/:B��=�ƻަNF��O�Rh�ez�E�M�ϻ,nbmuD�4P�W����[��udo2꽓m�_dm���5��X��̺��b�'B�|.'��c������/]����.��������E	�Z�BK��zF�}�&��+4�3%-`�	$ym���	��͒�̰����k�E��a1����(4�p����$�	����znu-�:w{�!t�^������:%�؅��L����UC���_bO�s���p�������	��	'c�Kl�ۮw��ܷCw�#�RO01��6iI�.ʱ��&�F����M��d���x:<�q���[;ItURC�����x��6�R����� ��D��h�^q؊\ۧ��H�z�W1� B>]eה+����1�{D�kk }��Ԛ����"�1�6g�
�!���{���g�H�-���d0��{�'+�p����53�i�߰�=�O��.Fn�ˏdC�Ae��\��(F1�T4=V���>C�̦at�W�S��H��O�̦�����R�s�,s���]V�f�cTD�OW��/��T!�n�8ym��%|u�v�Gd_a�[�1<�Rn8Th�D���ʻ��y�[R�x]���n�&H<Ő�|���ts�jV�tJئV �h�w����J�Z0ǖUF���Hٻgڷ�4][�92ve��1���g��i$mlSz��Og�l}�S]m�|ko�vlU������#Y�^$���!^͛�*�:�))��ʊm��-Z����ۍ?m����1.�C<��Υ���Js�Cv�^F6FP�s�_(N�RD��J�
�Gz
Qy�KG{��<�f�Ϯ;נn8���a|:qs.#�jy���?o#��=Wu'U�Ex@�e��r�(`���o��m���_����qĩN778d5�/k��6���6yւ%���gE��|O�����[�)�;v|^�^���kl�$迷-�<sM��~zF�����^i�x�
˄�^������C����aN�\r�%
^FL��',� �w��Q���I80�l�	�my����<k9�l���vh.�|���|nݣ�u���<kR]�;NjU�0�
�K	a%"��a�[�bo���W���
&�R6������8����#�F+�vb��7�q1\����FK|T�5�b�H1砇iI��>�����H.�~`��G�����{P�D�DlA�{�:@�Xs�k�s�&�ӧ"6K��R>�:��atR�V�ajw�3�`{�n%U�~����/j��zC�BV;����<�r+k���w�-�z+�=v���sf�í~O����"ʘxk�ad�
W��J��<y~W�9r$�Zz��-q#H撌-c39]��}�>���OM�x'ׇ�qJ�v��xJ��x���؄m��.u�qKwy=�*l^54>�\e�7�s׏AS�9�:'�b<oɩX:}�~yW���^�8�%�Dڸ�і��-
�=��1@��F7�d	EX]YyU���6ǐS�4�0nI��.6)�i��[Z�h����0�PyW��S�n��A1.�GpR��$������������(���X�v�l=rږo�:΁s�y����$�y�I�#�P���WCHA��W�J�]_w�V��	�vY���%�����KE6�N����7�x�s�RK�����F��%C_�P���'p^���%.=$"ٹ5������s$%��;A�1T�G	�$���������LBuxs��
��IP3Y�*!�W���S(����bXB3y�#$I
0Ec���"�%��������99e8���"��ķ�!ӻ�_�k�9�	z������O�w��u�f�7��xl�%P�w���hw;h�g�l���K�(�(d�*m��/��7�)�R�{�,��%��:�Ϯ���;��a�����[��� �Bñ�:=���~�w�	ޙ`��Y`B��Hf� 9�;��\��/�S��?�o����q�b�m]�B'��J���L=�`��[�7��cR;*��b���8	H�;%��+Ʋrh��H_�n�xջ�[�8����o�t^qܢ�W�8�;�A#���\Ȼ���ܫ֛I�+Ati��!i�C��ۗ.+�[(��	�*Bў�E�bg��_��T�h~5��Ҫ�^�_�=��Wb몭�*z��q|tG�۳Ň<!�L��:�o���;�H����>��f0�!�h�3!+����N0�������[T��$A����2��r����]py�H���Yy�����a��<~~rl�YA�4��Ћk�r�ߎɅGsQ��Lބ�<�ѫ�K�t��=GPi�� �m3r�^����H�z�^�3����u(�=cg�:��J�S���{�����c���-�m�E�w�<K��ĵ��h�~��#�	O"o�/9171�z�
���A�ή�&��[������B[߼�HS��ח���� �h�2�;z�������`@#�����A���/��ߎ�bW���HSw����}��}�����J͛�T*>!��ߘ����*M����B��Iy���p�躯e��������U�@��z�}k�n1D0�\����8$�Ol�0!�*�>u�]&#�6�w)�B�#��D�y{�3P��ͻ�iԩ���ILF�|a�#����]k�6���B
��C�)���_�b[4,��z�Ξ�����"[�c 3����p���B�����3
�1d�u��n4�5�,�V��u�9؉ 3మ`�v#Yɒ�v�����{�P"p�$�J\�D��������V�X��$g��Qp��0m���Ҿń��T$W���+�{�d�_
�Z[ȵT#E��v��RP���"�'C[��:��ٽp�ػ��A��SA�(��Omm��";�]��J!Q��n6,A^�Y{�O|@a��A�:��8���)߿���ѯJۈq�����w�TD��c�QS�}�&3`��O��
�Ӝ�"�i�6_}jL����&jQ K]�����샰�5�v�T�K��j�Y���g���
��`��r��g�j�1��`�vT�ABo���r������>k�}�6 ����T�ǺC>F)�R��
J'��SzE���=�'h�TD �^}=�o�&���4 {zG�w�]����!߆���Ͼ�'�&τB9=��,8	����T�M�Z�=�C��ň��B~3��Z.0OEE��#'t�r�γ?s����-X'��H��;�%�ْb�	KQ}�	"���<<��]��L\���!^�Q�Ar��
o��]��z�u_�{w�ap�� ?��$l=�'?T#�5@�C�����%?�Lbα ����EU�W&�U#���!� ���f
 /H>�����&]@I����5������{���A)��^� ��S�Dqz�6����:Т�Q"9|�\�n�M����k�^ۿ-�B��T"���i�wf���79:C��Cˈ���\�"e(��a���qɁ|%B�Sr�ݫ�C�Z(�����{,��,Q�T�]Q֥䄑2�8zF#_���Q�yyB���("��/����nR|Q�h<�8�(���:�ةϔ#���$�V>�y{���y� ��\	%�"�4s'�%�7����*:��{IrB^5tA��kj,e�� �A!��	��w[c��*�L�HC#�{�a�>���U�#k�3=�Rh��A�����;p��k���i�${��"�_~��4�؊�<��@'����o�:�x{m�22��-~�ar�;m�9C,��s��Y�m�1���X䷋+����I��sh�Ĺ�!=f��)B��P>B��;��C�#��B�D#Eg���	@�����:�?;5g���\E�E�x2'h��|6aM���{��gj ؂�7�+����@v��ΡL�=��4$P�D��Y�1a�PT�T>D�R9@8{)A�]i/��|�@��/a�E0�� ��k�Z�,]sz
ӫ�AE
Z���)�<�UkS����(��p^+��;��ɑ�F��\)7Bʠ�Tw^G�z���CL��B$�1[;c���L�XV(����D���Lj�r	{��hHo3�w$�&__�}/d�$yP9~Ud=Q��P��h@VBkՀ�ne���O�u�iX#���i֎b��Eq�E�yƩ�l��3(I�|n�Y�7�5C��A.Z����(�䅑�<x���Y�3�W���S�DN6D~�o��W��z��������Ev�*n����hTI�)+dr=짝,�PDDJ��/IU��	�L�E�n�o�MpYQ7*1 �k�R�~�Y�yB�0,�{$�^�l땃D�9Γ���������J�����~��７�Yg�oƚ	<3��8c�����H�Q� �@!TH	RH`P��6Ͻ��Y���ӝ�Ӌ��XQ��cF*hdE�q1UN]
D�pC��MH����2#�$�(�, B��(�w�2 �;�0�N��D������;  $�Y���R@B_�1	@�h�d��IU% I@�q�d�� �(B)�\r�"§�b+��+*E(��L�JB�i/#�J�#�@0@�H@�dR�?z�Јv����h8z�@_5�q�T�?�SB���/P�.����/��1`FG	U�C��[�H� �O�BRЎ��'�~?q��������(����{�O���� ���AM
q��l/�}r|�~�`�y�}D*���O�}����}��������~#���{������ߣ�?9���������xh�zI A��?��Á�U��8���_Ͽ�=G�s��������o�����o�w���տ����9�O���z�_���o���4��a���O�C�x��_��'������Wy�s���S�g�	�_��?��?�G���?�9_��TP �����E�s��T+�!��1��׳��o�&g�o��k��<O����@?�i�+��������y�f1�I�|��)���/߄Ic.e�-k��J*�욻��� �����������������Q�;��)���_�Y��E�����0�ʈ����2����� ���~Ҥ��G�����Ê�j�y� ��`�PgKr Q�e5)��f����~,��9����1�����n��Ԭ�d���D�a���f&���#�p����g!%�93�s@�V ����@��O��1����b߹��֚��q/�����f`��k��E�����Ě~���+�^���f��=܇~L�$SD�@��3	�Qy�$���Z��m��4�Ee��퍙u��=����t[	A�P��X�C�b��o�'�����o�������������������@��R���I��|�����0���<"?�ß���ԇ�j��D�)�J1����$��Ј���2kp�w���	�������&���$�����%8 ��S��$��K	P��-_�+��W����dx����d�Tޣ~n`!���3��wh�46OE
o!;ª�Vy�-S�����+�?z���E7P�O�q!Q���̽B�2�XI�L<��\��T��A�a���DSQ�� G4��=��5L;#�{���οO�{�8�� �~>L��u��`�J��_��ݐE?���_��_������/����" (|�{��� �!(
a��ۖ.�����Z�4�nr��h���IE3XV���S��G�)L� ������6��E���|G2�U��I���:?v�"�ħ[�^�  �IZ�Fi��gN���wG�B�R- R��p��e��׻��ۮ��ֽۜ-��`���2�qA!��6��l��C��L�]�.:��$Nz���y^w+�tb�+�+n�:tswv����]�E��"$����	/Y԰ug��aS�y�Qm�4��3�/B��8�C��d�[K"�3����YlX�c���j4� ��q�D�n��W�b�o��S AR�A�⪠�<ۛq�T֖,ԅ~���������(��˥I��|�9t�����)����li<8�O�Q�o6�j�<�g�t����qm�E�Ŀ�'��k@n�a���{�P�\C�g B ;�dp�`� D*�"�{���Zf �z#��ה!y�>m�DY0TP���t�x���fXi�Fl�ю�.�)�L�� ��$�(��) �<r����kEp�&a�j�Qj�8���5��]7_Khp�x�	4JHO��q���~8�M'߉�@�&��|��6L���Xm;qÆ��dr��&F�ǖĲC~����np!�,9n�$�Mc��I�����Y^�� �ݭr�""*�d��נ�VbgUMcӣV9�ji�їn#�I\��-U�Q�X���cE GI�S��>Nl޴9�
h�6t[�4�x<�QP;�QN�+B(P@��Чo��2����x���&�p��� �ږ6�,[�(�Ӛ�Ѯ\����4_����k�
�0(��ޘ�b���2�$Qz`�H$��B!` !T %B	�N9�S;�RSM-*d!��(���}��g�����rš0cE������*�t���q��C����x�N� 0�n¨R(������w�{��D@����(��l���DiD�=�����\�C������ki��=o�7�/����;��,�����C��O?�_T��J���J�����k> <_�8?s�}׾�<M�h3����ߝ�n�Pъy�gn[���T�cpt��?��"����Ϯ6E�oM��6UHJ<�C�Cc�QH8�x:����=_X���������K�z�/2�Hx�'0��������y�
�N�DT�v8�0$~�྅׏()����xh_��?����e?�?W�8��,�)��C�	�E �r Gߏ�y��N�י���?! 4v����s�T�$N���J�y��� �W?���ɿ�����h������<�v��{�}Pn�����?�@� <�
n��т��n��|w^���I�;�W���O����/��0���?���Hw��]��)� ����sO��σ�䠋���<}a��m������>�q?��z����=�����Y
��!&*�>mi�i��d"��m���Om�����[FF�&-�5kw܉)�`���qT�'Ϲ���c��~y�6Vu!�TDDb=�(�'!9� ���0��C6�C�Ȉ�(��+��`$��H� ���: �)�I�2������kF�϶�ͫm���mg�5e�;�9� ��!i����
�"��(����� ������3���޴ �����G���QWר���� ���E68wh��������P��?�ݟ㞭 uw}��F
s���  ^s����"��0t�t� �ࠏH=H�Q��~]�߈%s��f����� ��5��֫d��X�& ��d-Ll�j0�
�
���u�!9}��ׄ� ��p�|1Ԇ���p'>+���8����(�⊰�N��J�=����<�"����LE2�A�����I/��h�Ҩi<DXQN�N��=c��kp)O7�ޣ�P vS� =�<�|�P�"� �{g���;Cz1N���9'��^�C�$ YxzM)�~��%@�|�1�!ޛ��C��Z�V�c3[l÷����t�~�0��;�d��T7�.u�N�� }"���G�o����*!ԟ��o��7C�h"dЏ���������>���2�⒜�����9*�v@:_I��J*�O��/-^OJxw}x�k0ʱ��/�.��wT�nnn-���W7w]+��6Mg9(�ۢ0�
������U.�4���y|�f�l� �"����J�˨��JJ"��֏,AO T;:T�ҩ�*�G�SnO��Р��쉡�8p�Ù>;�AEz+�:P�v0�g����@���ݳ[)�	� 6�Q!�S�}��h�GէJt�@�<UV>�xV�s#Ϊ�1gH���w������x+��}o��4<�䜳�4a�;I�Ԩ�n<�֮Q9`�%?�����}��' ^��P�T9�K��A��*`M�u?���<TA�мD�'�L8hSS���I����HB���n%�g�!������K��ڡ�j"�|���S� ل=�ڏÁ����`HPzc���8�y@� ���w�`�c�5���
�!�vߊ~?�_��7;þ��Q�T�P��H��v�"�zoB����5����5z�>H��!�
p�B�M ���ET �x"��Н�+�aP�P ]Ӳ(���x�w��� sʒ~+�<��qS�BA��E�:��v�6aߠ!8��t��=�}�9�q�sl,��Fw�kCո�y'B���m�}�Pu��;/'��;Z:3�:�h�s,��=�9ǤܐC[�t�� �S��Q^`4�>/2x���<A��;����W��� O O,x v i@d�*�=��H�?Gl:���w`s�ޝ�x>1ވ)"��қ�� wP'?y�������e�0��@��<���^E��+�)�?y�'��G�4��;��I������ ��潶���v~���S�;=��"����<��}�����^��H���_����tq=����m���^����¢�����/�� "� ��(��2"����4=��/�o��#y�OxX�������0�7����P���'>���Vu��"�|pLT�X�`��?��O����~����|�?��hO��'�?�~��o��������h���_����f~��>��{�e�o����_�/���~K��o�G�~Ͼ�/�'��~�[��]�=�������O���~׏+6Ϳ7�{lۏ����Ϸ9�� +��iװv?��yq������d9��Z~4?�$c���c��i	�����[
�u$�q��}��f6U�E_�R��_�c�8(>G�<�C���]*]>7j�|wpp?)a �

v��&!��%��h�� ���U��8w���k�`����>H�ll���4�,+� K�0�>��7�����I��@��φ|b_�}*���������� �?�b?�����,̶E�g�q9~�a�7���`��׳~$j'�ۿ�/���>`�|'������S- ��+�K���_�@�����{���I�}*`�
 �u��j"�4
��f"�Ӟqӡ�&Ȅ�B��*��k�-��lZ7@�U����\6Ӻ��v�k�}�<�x����|_�|��~�.M
$�H�
��
�,(H�(�|�����s�G��;�3?������w^����
����>w����;�_��]�N� ����8s����{���u��!� J�!  �$ @��, �� ��7��&��	�����u������N�w���_��W�\!��pC���� ��������������g��%'����+�� T���zŁ����|���b������:`BC}�9/������ 	�"@�� ��Ȍ� ���J0� !���KH&�dP��<��0�'�����y������9��_����N�܊�]B �W����5�^>٪���j����yG����}��ήnc�3���i���׋y΃�zN^G�<�z���%ߠҸ9?�������O����%{|�I._g��A�-T�9�h�F�~kI���>	1����[膈�nj�75f�Wb��j*d�0)] +*���+G�O�?���6��+ޏ�H�6�5d ��s������Qb��x��BI�Bj�\��5��O{\T	�V����D��S�w�fj���=�Y��P��!����
��O����YFu���P�S)�D�1�e�t��Rtci�����y�����Lwb���>��w�g���/�6�'1�C�z���ݸ�\u�B��eԈ�Յ%���ʓ�ɩ�6���ΐ��v�C�a R�@d P�`88� �����Oޒ|����$�+Y�2ץli����b1i�^�i�渃�n���#����o\�ز�F���2��*�/��¶)Zɮ��Ɵx^�Z�9�Kb�O��c�+�?�s����Q����X�����1b�9��`��z�p��.LYό� �e��,��F"��^U�o7@V�����Ci���'���-R����P�I��_�j�;�O����=x�G�u�h,���<@,����[<�Z�����3���m�r��i�4i��- s��z�;��q���}�{/�YN�h����Fկ�T�AJ?��q�s��M$ћfr�6�Hg[��y��|E�sX�I������9U�$�I�ц���f��V��&	εc���F�Y�[l�:�7a�*nmMUЕl���ؒ������8�$���8Cs�6���J����S���r���S�ﵮ6�c�0�Q�9��I�u���hI�mbqij"q8?��?��R�0��|����e��P,�y
��:�F������y΋%��m�b�+�n�5&����.F�3=opv���6$�ޚkj����Z�Ԡ9��"��n�����C}�x��D�e�6|�\�L�Eΰs�?����O��v�S8�Q��!����Z�~6��Q3L����A��dg���5;�hՙ{?���O��)���;���'Ч���$5u��o�����F��R|7�㥌�:^��Qu��!�g<�xϛ6�x��=q��~_Hq.���Gx���k�Λ������
�Z�M!^�Ԅxt�+j�-^e��C��23K��:���?�#���f1�y�^Ы/���;�E�(ݫoG~8���yl{���lT��Ͼp��Y?m��e�$۶5�����_=���ǇȿO�g����5���k���5X��=��޽x�w�������	��l#om����K�j�9X�l�P�.��-p/����v�2leFb;p���;>o�*z����>u�n1�`$˝(��ꓣ]F��Ԗ��i_�m�Xo�	�������ng�w�;��N������8(s��I'}�~Qw2�-M� �\Y�j,��4m MZ嘤��]�f��mh��&��Vy�Lö `p����ow�~��o~���}���Tէ[��N��v���U�>���_O]����9��������O(��߿y�8�Y>�#�?��_M��<���9�S�d�{g�ꋆ��}��Q�;���`�'�4I�^a1��/	Y;��B�m~�h|��;y}��<c�|7y�q�Ϟ��k�F����Wʹ�np���D�M��#OhN��*��'�J~�m0���H�F�Ҵ�T�+����;�7����_<{o$��-U?�q�\������z���kK�>�5M���?��:�q������N~~s�������G�u�T|��8��C��q�=w�w�Ϟm�n�>��VDk���a�e[{�A�m:�:�(�:�K�ۯ�G�F�\%%Q4��x�d��>��≨l-/����)]�^��Z�o��s�n��\>s�٤��n,ժu�"�m�y{����~ޤi���A��5;R���%���~��$��uz��ZU�уy�����çl��j�~0�c}>�y�%f{���s4g�ʵ�7�|�n�:�m����adx��������GA�� �hl��h�F6�D�d����@=�H���!	�	 �aFE�VeH�C�]�]��R���A�ECx��-�ݕeX�V�C,%�}�-�c���^?�){G�GV�����J[��ߺ��{_>��z;|�)��Q����+/����I��������/����ɽ��o���_�������R���������>��/�G3�V���o���~�$|�i|��O�z���s���|s�z�վ~&�2�$}��m����e���B^a_~�o|�Զ��l��'�<��[^}�6#�������w=v�����~�=~>��^�z������K�.���U���d=�;���"ߏ_>��ǐ��������Y��~��{�b��kl���緿n��o2��z�O|�lS�Oo��^���+�-���7�������R?=4�rx�ϯ+o�Z{��ۼ�ڟ\�'�<t���=��xOj��ǆ����7��|<���ߎ�;g��h�m��<B��1:�[�����to��^e�=���W���9{{��S�^���r��-w���ח��L���(�ɚa��<�rLC�Js��O�����_�o��f�v�����_�]-�������pp������v2�>��Qp�ZƓ���d��#*��1Ѵ�Lƣ���)�!�B�4[-ۥ��r0�FЙK�&�S�3Q����,bB�?����;������^��o�����~�HÔ;F8�oL�h�I.в����@��ü錦�axƖ�J<A�`H�!�[h�h5�Y�|�#*RD��f24\أ@P�(<m��ߏ�ֿ�W�w��7��O��Ϣmݻ�����<|�k����������ޥ{_��������_��c[�X|ռ��]��Q�n��~����XM�6�A���=�82ǣH��cю�$7�_Gg����q�-��0���o�/�~Tǯl}\,SR<p?��p�!�62�ah��/�$i�P��e�Sa������~XG���OSť�Q����ߞ���\��=|���_�_[z�.�6g���r��:�Wǟ��^�!eo�~~s�M�?]�����wλt���n|v����R��Gm�{Ϯ�L��(���7I,*�ю\
��M� �`LRz�����9���s���G�U�x�?0��T��1�����ߍ����'���^?4�R�������ժ�'>���=������}����h���-9��_��y�-􃿮Щ��}����?~~�[S��G�~ʕ��������=s��쫝���Y���>�~�:����|�ә|w��S��M�oS���p>c�}eÀ�Odaz�&A�u���hs�3�0G�1X�i���	�JJeD�$C1&���Q�!�NY�bhV�,�ͭ��}_����M����*���3
����n�ۯo\|�(Kt��S�BP,�q��q�}�8)XzXc!���LO�!�F+2����,
�B*sK��
�<� x�zv,�!qfL��1�E6g	I�K0�%,P@ ��њATTq�����F䆍1�4Q�Ϙ�1�ASH�K��
1� ��&y��˭4�I�������33������"�M.2�#8(��%$D�`���k�:�@�2�bUhx�*"<�	!]u�%�_i�N&OdOJw
%@H��"K&�/	(�����ꅎ�K{�)�B���68�H�`x숐�(*a4˨��bE��}��9��[����h_���{v���՝�������~��PX1]tɝ�'��fR˄#�����҈��!�Œt�U3��ѐVEU�L�S`H�ã
�E��h3�Y���L���F�s� �0<�>�".�i&ErRKg�.4Q��$w�zr�"s$-)�� `N@!�@�vC`"�`�ܝB^B$f�~h�`!܁tM*C�Mf��� ��qvb!�Ӂ4_�)cew
	uZHƘA1
�������,��sn$|�N<�;��|�9�G���2��+$Úln��P�"!+,��j��b<���pe ��,D�Zr��O,K %�T���&
X�� !�q��?�|0 ||���Hn.���P&�T2Tj6�!.�����nfQ�3Mqٛ&��TipI�X;�T��|�^�+I�r��pَ �����8C:�O�)p�uc�T��lx��G�%I�nZ�4E�&��)�NyeS�%�bI�1�@�� �+d��(��{΄$�*��|�� 	�#�M�J}�5^}�*
�J8�6hq^ASTV�2�P�݀�`D*���`dRMY��f:k���@,2N�F�\#�x�1�d@�D%�%�f*	�5c_-�!�w�nT�H��LH�%Z�LP����R�cЮTH��U:��5A�V�WP��Y�����oTp��5�v�=`Q%Sd"�a����H�Na�Uԕ�%���*Y�3	�Mm�D*�E�iRB��h�P��F�+R�G�\$�X�T}h6"�R)2�'�!�+T�;�(���2 �"���zP@uc�ǳK�:�|J��VeA�y�COZ�G2F�4�rH�d���C��C�,}T�h�6TU�>�i(lQ
3��HT�3��MM�е�K	�LJ/C0#�9�A�ilscV�I��XR`@Ƙ�H�,��9���T0�����s������El���c��Zm�	��<��jc(��8�A#� p�#CpcK�(�uAg�P6G6J�r�6�k�A�t�����6S�` 3���mV��FPY���R�j5H�I-e]4MZ.Q5�)@P�Er�btʪ9�U�݉'� �] A9�H�4ڐ��#��.*d<(��1���%�4�ju�>d*�LT���XI�Qg��Om�Q>�	F0�S�Q4R0�K�#�\�k�q�*%�2VI�^j% 5	�H��h�$�͆�Z���Xi(	D�˵@g6�A� W�  
B$ B�@#*B+(��H�#(ʰ��B��"���_����Wu�����ϯ5���Z��S�3�zT�Pj �d#\��U�J:L�.�0He�)h�8G52�.hd���@D��T*��.�����0��n���aI�.�"���!��Q�Ij�C�kG�qȫT#|��DJ�I�TX�]�LM��ܡ�3�.UAw�0U�֠i�=k�"ժVR1&u���@Fa����r�r�4��6$������l6��@k�dd��o$�D*�]NUIf�̂�=;� ��2Z|	�s��T¶�HY�0��Jp��e&Q�I�Gh���U�&�{frCT�ŸfF9J��nՏ.�E���F�[.�R�B��,"�)Ol���Bs�%[�#)%q����S�M33AkAuw?en&U\�#�N�͏������
�+���TD ��V��[�4�N<QGJ!���iC؜�ᵉ�5�®��-����4aV�u�eNL�v��qUm!��d�4IL�@���Cq��.-T-q%	q2=���L��3P�lR%5��#N�$Zg_e�ky��<Sgl���bb{A�9M�h�C�4�H3y����DCH�Em��2$k���(/N��:�(p��I�'9��F�a�SY�/Ub)Z3V^I�&�ڀ��b�Φ�`6�o,[�����L#�V�@DK:�T��D�W�l%	4/�ͅ�i��"]Z0�5֩v4��N<o��
)����j�SBQX�?DЊ�cl45T�(B/jR�vBRԌa�� �㦹O�)F!���eb 锉X`ǮA&�aD�[�Y2�B��S�OI�H�H�A��OQT���D@[��J$D�E���CҾz�^���:�Z���".�Ώ)�>1ډ�����ux��D��E>�Y�J&j��ZH���E�����Q,���R��J����XzKXی�h���]�����u������2��R1�=#�+��l�$�@���d[����Kߦ	��B�z1p�(�'Me�X$PDaE��R��A�D̉��vw-L�G�a��H�j�"X`.��~�K����^iEUqV���8	s��M�&�%ƓQ�8%��p��,C��R�v �觝/�+9�M�R�C�MΕ��d��������a`n6�k���@B �bq"�c �/A�I0K$��Q�`�T�$�F4|�z�ڤ1L�fV6�-�Z�Xj9fr��Ρe�����c2V��r�rk,����a�:�T���	S�:d�UkÕO7C����$���<�@]��a내hm,��̺�">X�Q�+��.�C�q9E����;S0�c��ȶ�)h!X)@"�".�c���� x��yN2��O�5@)�U�Ɖ�!���4Ēr������I��Q��L[�@a ��[��W��ԩ2k��j��{��IB&B�pՃ�5�P�zAUt#��HYX�+��/�f�ڙ��̑���i�h�T��)�J�즊� e��$2�����!����d_E�Z�q�%9�14Є�Z�b�%��ʗA����	]��
��5`�gP@�/�봔EI�H�\]���m��N �R�pʨa3�Di��0&�EI��5z��I�9��6�i�`��7K,�d��h�Bx*����PL���$���Ř��D������H�R��rh�	&��+���B��1`�U��,��/	�b�m��q�)��;�2��\��>w[>#j �h�C�~k��{���F��%b�>	I*ɹ�ٱ�^2&Q{5Q���-E�E��f�����P��C�G!А1C��ϭH��1�Z �Eep��Oa&�[s���<ݏ
��$��є�� i	D?(�a}��(��K�9R)���$:8�{$M���jj�xh.Ԡ����M���q�80Ĵ���pAy	q�]��qbj�f!.�t�@�y���fv�Z�h�]��>?� � ||  ����<eg�L��INN,�d�o�(�fR��i	,��(v8�P�bh�� �UYT��l��L��l��K��^+�=���[�5fČ���t�s���3Jmr�{4H��/�:�;i�O&���<Z�E)/�Ճ�+��g�b�mXeɠJ�:Ew��K �8�50�%$
�/�6��ctO鍘������i�0����Ԉ�僊ŗ��F �q��<��zÖ��54���;o٦m{2@�4#*�"�_:q�-+�i�+� -w85M=�;%�k��4zd$��~�Ja�Ms� ��$VA ���5�o���dk�"q�U���dN�y��t�3��;4��&��2l�Ȉ��T@�(S�Q�����+pX���ĜF"�sa�V܀���$� ��P
a�7fA�t:�� �v,�G�}c�)��)X�kAQVA�:��v�HS��ĉ��7 ׆��5�p�%9T4�]2	���Y���F	,V�4N<�N�6,s����\DTV �;&�c�<��� �A�@�e�gX� �b�Qɫg��{�A�ֺ�i�Z�QҎH�����I���e7�ha�p�6��N�d�cH�E�w,V�7h�,��e��se�<�]��P�sJ��+R:�r�����QU�0���9$JsKd�5�L'tt2)��B���Q*��cI^m,bڄCg3a4��U�c���֬Q�M�F��\��X�n���d]m21�R�iA*�V�,0�gc ����Ly���=w�{A�0�:dF�QGO��5���+3㙝wY+d�yd;��i��S�i4P�Zk��.�`L��gv��T��f1�h�f��b�Ѩ��э	`��.>�.g��iҺ3��ہ���~�̑�{���!ܺ�n�P�h�5B�U��{"Y���n�a���adR�qn��^��F�W��sE.b�o�b����I9Z;�R?�z��	<�\�R�`�ݞG@�׉D�$���!����xl<�2kmd��4��뷩@���r�e���
�XΙ/��/#�?9����D�Y����$cpȉ��@XC�\k��tbT�(�A��8}ge��`�r�̭�,0����1u~� �?� _ +"P~[���.�([@��H��ė#b�� ""��N�3�K� ���U%�+��0�a΂�T�`��־�9ul���iR4(VKF�n[F6��Ȩ��\����*�\���kr���~�����g��辣�_���ـ
����A�lQV�kY��Z���*��E��h���`�V��X�12�4�E"L��� (%"��J
�J�R((SCB�#B�H*��dը���X��[b�E�m���F�ѭ`�V�U�[FմB�@���J �R
%"
H�P)@
Д��H%")@�H+J�@% �J�+H)H*)@�HH��-�J�%(�҃B  *P��E	��rhD�MB���M��"P�%4T'x�� �E��	A�B~x'�����N��������;~������>��{�~?�����������_3�~��}��g��7����}����ξ}U�C�ȸ�E��3S!A�2��h�X�e��L�&�4�))b$&�IQ��(I,��Dh� ̤��$�����i�%�c�L`lAS"�	 �HQ@H�""A%4�H����&IaB	�"�d�M11d���$�M���3AQ����d�@d��ʄ�.�!�C��H)Bz�2D��#�r<Px�Y���o^�������>���
�� l �C�=T���m :�5#@����JPd�8��j@CD)R�P-�2�R)�(��gdA� ��d $�m�
rGP+���&�Du.�PaD�X	�"��� 0� �i�Vw�@!��T,, H�bT�	��A���������U\�$�I(��)�@0�FF���k4H��X�@�!e��g&���Qh%'F*�Ty6��iX@�@�N��U���������?��m�^���ð���#�~����Ǹ�>c���xg�9�����n�3�}'��^���g��P0W��o�7��K�E4�쾾�(QD����������p�G�������w��c1z��C ^ulqV͟��$���i�sTV/��_��������T-���D�?�t��I�����;�+��l����qa[m�����d�Av#�RA��sG�<ކ��;�y�Z�J����EF9�+��a�fQܖ����Xʨ(X�AN�Z�Jm��P4�X h4���i� ����L��}���(�c׀��§�	�Y2n�,:GJ��ks?SCI"+�ޒ#i���ڝ1�����|����1�}��oc-�*%�6l&�+�xs8K�݄�"&VU� K��&���z϶����V���L3�5��r�v�\�n�O����X�1/��8OD
̂�V) p�u����H�e��������2Gzm��
ۤ<�pk}��T��R��C���@|g���u<Z%5��Ǚy�ATF�,
o"��m��\��}������?n�h�>���-|�?1��gl!dA�ؠ�BG&>��%��֑Ie;��`f�%@UV'�Q@�Om������ ���u�����j��NO�P�?���4l۶keSD>���J����˭\s6�eϣᇃ�
[v]���n��A�Ŵx�r��������n��\d����
vAh�rG	�=�E��n��R�"E���z+�5h.1t)���.G�Zϩ7��4:`?sB�� X��ݾ����.�~����vMGWԄ`��b��dm�q�
�f�>�U�d�(~`�a/[Ӫ�^�{y���b4e���V�)����V?�.z��3�k�F�t��ro�H�Ee��f����]
��;�òc>��G��Mږ�6�"���CW5c<[��j"���� Ri<Gj|<u�PE��#z�Gg��&:��W��M�\��*�0�^�ҤA���ad���D]q�g;3�٘Z��a�֡�+�y��q��vAǲ�T�oݥ�\�ׂ�İuw�v�-�
�X��n����GN��]�8��<���nvDB���4 ��Noo3:v��%q
@k���"�:��v	^M!U؇�cm�W�6��#f�=����aYR7D�@+:��p����n+:Q�X����M�E&� ����������,F���3(��5�b4Aw�$��V:�?�]F9U��8Sn3�`ŽUR��>>����&�D��4g��1ڝe�A�U;������!�*�������>/X����������?k�J��Z��_=��:�t�.W��`����a(��*�*"� 9"��R����9( �EP�S�e2�U2�T�Tu ��� G˕T<���zxUT�:d@�EC�B&�#�
��Ż��r�;:�m��U���X��<��|o��}�}ɿ����G���d['f��Г-#@� ���� �a<��fB):0rl���,<�{?R.�|D`ZLXM5S4� \�D��9)���+�ˊQ�5�W6��|6�{{�vC��;�@��%G�+���ɑ�U5*�P=J8�i�D��b��L����.x������������������������������������>�E/�R��w{�{�]�ZVU�z{B�@  �Z����       O                �                 �R�       �J���*��l6            FR` k@ (vaf @   4�� �    z(S���=     4 P  �z��    �����   �
 �r�   �B��    �DR�_  .    �Ȧ��   �    ���.    �<                                            �}      ��    �o������l t � 4�MD�	"� UE  
  � 
 � 45���J�����(*����T  q�@�� > ���k
�356��e+w��<�KP	) n0  IJr��@ 4 4 4   =�@�}�#'� �    tR�>��t P���*�� B� h7X �     '�u� @     @*��     �)&���	�m ɩ�22L��M�Q�)�jo)����j'�����ޓқP��<����L�4� 	�� ��)=@=L�P���Pئ�G��ɧ�� ё�hڍ=M 4�4h �h�������� ����R�H"F�H � i� �        @         �@  O$J��"�� �m������4i�� h2h   F�!�@i�F�21 4 h  '�R$��'�)�Tz��6��OFP����F	�CM   L&�� 4��h��ѣ�  4 "I@ &#&F�0	�&F�0�&LLLFM&�����M0����I�#@�?& i0F�O�1�t��DH��B�F1�q�����.Ma���S!m�J����)�M�6�-X� ���[,��`I�i����id�x�7z�2�ӌ}���n���̝�������]ץ6;%d�3we->;s6�Y�J�8/l�y���$`A)���X$H�u
>�Tw_�^׭���q�c)t�&�F$��i�N]��k���,F̴(+��NbBf̀6%�	WU��Q� �5ǜ��⍠�����[`F"���A0/uɮPd�Zh�f��9�DA���0+0���r�HDH���qb:Y�MY)V.(��Y����)�ě���_�6L�>�I�"(!��!�C��\l�u��*ҭ*�=y�Q]^�	V�5������V������ ��f���;	�x��O[/��g÷�����9�_%䨺D.�E���� ���1�l��Mj����\�inJ�"��I����1�=���Va>fAL�PH+ �	�$�
�&f���O����c��R6�~���}|(n��7��>�e`a>��*g���W36뛓++!u������1_��!b�
�ᐔ��2L|Ꙭ�?��|�*Ϟl2&<��슱U
 ����'��q1N>߀Y%��s��1k��B�vt��Cՙ`�&}�z��yo��=6�n}9�33>Y+,��ɒd/��+%Hd���!��p��&������� JRzX�^Q�=�BwV��ަ���O��>Wɢ@�F��(�<*MT)�=+ޕB#?�[�ݪ��L�t���am4S9��=�B���Gy�M��'�$��RbDL�d�L�Ab�Xp�B��[�24eܙ����K�� �H � '�����^3�w�"\a ��!O���|=���P]�#�(�(��1�Z��"up%�w:f}T:t�'�0�͟�P� �̿M��6�i�>����bQ3��
�b@��%���C"E��B��@Q`-e��0��`Eq9�!yDAr(��!1DEӒ�̆M��l���5"�!�#RVE,�2��C�_�������2���BP=�jJ"h����c�e$��l��������D����1)6��fD=����4M�J�=0R�I	ad{�[��|4�Î3�d+�l4	���~�f�0~�ߧ����tWƩ!J$3��G���4���K�0�o�I��{ɬ�Ak�Bʒ�#�������$�+�,��tgs�	0d{��\<>��zK�����̨s��OC:������F�Ŀ���f~Z��L��0��pR'wˤ���'��s2s85�R��,0��|w� 3s#�P ��ӽ�����&d&�!�f�,����ʫ�u1a��T$	!��[%V�Q�b���?���#&)qD@
YfdA�S��P��R!}�Y�K_VK�Ć%���Kf���fa'����b�S���t���n�%����?t 98��N�����e����ހ�z����x/��n� 
��>-���E�e٦�㉺�M�e���#�Qӳi��6�t�ݞ�wsC8��8͡e�e���hdB2t�d��8�$�C� 6wL�͓7�F,�;�#%���fN�cɤ�c� f�V���� H��h��IHd ��!	M�ޅ�Ze�M`K�u���!)'^����[��=;nt	��6y��@�K��Ȯ�v�^wd��r/Ѣh��.rS�e�r�K�Jwnn�o7�'��]f���r�3����蒐͐z�s>�칒��/��Ѻ�vuZ雡�΂Ni��g���}ۖ@ @y��n��+ik�ĒL��	m�9�x�r$i-w�� �@�U�� :��h�	�9�i����F&@���!X�8	�e�nh�8���N���*đm��X"�,D�.��t���2�r�ð�0 \�у��XA��
D�-��6�`BQ
��J�ՅN7P�vX��vk�ܔ ct��rׇ�4h��5!L��$�w�aĬk��"�k�íer�ި����1x�7j&�+���
Ga:��%'2�i��z75��;d�nUi�x��d�GJlw�HYj�	��5ٳd�gCY)H;x��ړ��
C [J��%6�cM���]���R$�9ݝf�{�x禒���;��vp��.����xJV�D�W��H1��n�s���L��6;s7�7����]kK�$-v
�Hq��H�!�D܈�
�E!�^5.��k���Mb��h�k���d@c	9��m�m0�$$RD�\4�N���"I�
&g=����ܨ �@��R��M���iE�+4�+�  ��TB*�",T�B	�T�Mk5��V�e�����@�����^�����ƪ���W����B���݇�@ Gc���� M���g� 4�@QF �F*��55����[cKl����	�M�^y���y�i��{� ��.6�f� �M)aSk��[&�W�ԤO5�k��?��s���f�����ß�3wǿ������w�{�1�/�{���f��#���j���G���D{Oe�M��?G���\g¯�Oc�,}/���K�l(��������k�{Ӈ��}ߩg�{Oq9��ߌ���=N=��7�?�y͟1�r�����������g�8�_���|�t�S5@�*@OB���|p���E�؀�w���q<�����6��{�v�>����k�?��?_?��0/�|�}�P��N�A�0���������G���/�B?ɟ�w����oV�8�3)�͸Q������~���j������G�G����݇��}�M]wC��#o��OK�VӇ���A���r��k�������n/&o1�n'[���!�(D����	 � (H"(���.���VS�@�z=e���_@�u\~�3����N5b�k=V��~�C"���Ʀj�M�"'D/��W�	�t6}�o�E�D��&~nW��6c��ӂ�a�MF�'��l��%��v��r"�����wa�S�����^�r� 5� =|�p�~xӎ �����;�	O���U�u�z� D��e@�#��Q�5�ǧ��_>_4��wSźE���7�ߤ��I��!��[}�]�D@����=c����q_�WC���"j�B��'>��_!���*u���� ��k�[�����;}!)N,vhN5���>7�m��C��7��� ���Y������> �<���[��p�M|�DDD��R��<z�6��'��>�4�esͿ������~�_7�;a���2p������ @   :w5��kN��PTi8-��9	6n�g� :KR%ƺ��5��]g��=o�<n��	X�)����m��bq�� �ן(xp�>�")�  }�R�<{\:�6��>��?��]���z��|,���� �m������>cֻx��� ��N�����};?�>�ޖZxtc��ƨ� ����[���+��������?���i;�@����ko˯�A�G����m��^W�|�_���cw��}
  }3�?�����㭓~���:��p�"'rC�+۽:���\n�=}��_Iwε|5.1ٞX|n���� ��*����}a����� /;ƃ�ڧ�b�+F>�b��/[~{��D]=�^�������J���y��{�����վy� 45�����Q��d�=���H¿��Fx�-_�OgF�ߦ� AZ�?_�����֘�Y�������v�P~��hokʎ���pߢ � ���~�6���mK�Ѷ�����m�����(�� @��_���}5��o��Rf�i��T  ����p��i��/��;?0-�(�WO�����  �c��͹��5�v�m���GqN��?�>��E�m ��/���Zro���b(�k>L���P� �xlAoo7^3�o�ӧ��z���_���	�}j��.����K����FkC��������d���8��>�m�ۢ D	�&��:��7��N2���B^>���Pxzx����D n"Ҟ{�����y�9�`�|o�x��O��@�4P����v�O�Ɵ�m�>���{�[<���6���?�(�Zϳ��������2���巚  Ila�1E��=����Ϸ��  �i�^?=wɧث�Gw����_,�d@� �l��*F��q�Z�W�S���� ���ɣ��Ⱦ<��xw��=�,�Ǉ�����
�\�_�h6ش���[���ҕ_��m��%8(����t}ayiD�����ד� 	������5�j21�W�����֔�Q6�Jl 3�ƣp�`�0%e�%Z�""�έ�~�^�3�� �W�Ѻ����n� �v�f�˽��;,�����K�/����k�:�0ڇ����7�����xux����3|�_ [^�[�@��e�f�xZ�+?�}v�"�f�B���~�� � D@7��ѣ�����J&]۬�0疓��l���*����2��δ���|]A�����"  j,��������M����<����(��4�Vĵ@ z�D��"��qn��)�K�ݣ�������Gy��G��� �/�I��zUD��!���bp�Xĳ�Q�oo7���Z�Wy:��OP� _��������f��++ @��V��owx����/�j!�ʈ���v���M����uǫy~W��{��{�����?�ڲ�~~��:�s�m܆7�۟Cl� <��ax=�jk�my��!��5�}>ٰ� ��S#�"a�m�q8��-�v���fn>��>�?� @��� O[i�y.�i��?~ ��ŋB�gw����_9����Ȁ� ����Z���l2���03T@�Xb�8�d�|ۭb�ˬH�Z S%S�͎��" �˻��v���&���am��wt�V����m��٬�T�%�k�z����̓�v�;X��e픸 i,	�D�H
�zI7ŷX%�e&𰠌��=mRu�Je�� 6�o���f�-�/<t3�a酪�w1w���V���I;wg�*`��4��=��1g�x�gE���aa�ɑ�3IFv��B_n�gfLr�p΄�7\v�[�%p��W&���A�ur��FT�ɮotnԒ�۔ ��e�яt�f��n��wGT7�4�l�7Y����n'��l��;�l7��!�9��f��RYn�74@��,�����6��O��2i�m�"B�I,�O�0m�C!HMP]��۳!���Җ�ź�&�h��ݵ`���*�aS�JNk�BD�/@@��B0`"�#"B���
0α����Ji(��a"�-��� k�^&��׭7T۷��˴����]X�ᵮ:bJ3m�l��wf���B�ܱ�f�f���#*��M�^;���̹ٶ���Ԍt��2� B�ApbB�i7u�z� �!�
��ǎ�d
�H-\�CIe�Kc �YL�,��7l��[gگ ��唖�a�����q�Z+t� I�	����e�!���;]��,F'�l-��<�7�t�ք�0�A��M%�F2$7�ŉn=S��PX��#��B ��W'm�`N��c�l�9�rNK�.K�u^*I���:��Z� 0 1X*$�l�h���dLQ����#9h�[	�Eq��k��9��Y4�dx-ʓr����B�L��aJX�QƜXa�٭,&�#)�����K���)��u���$*WDu�[�͠@|��H���l�f����,D�P��%��%�l���i�-�N��������D�l�b���e1r:���6�n[�.�9Dx�%�V�f�Wltp'��i�� @�sKݻe ���z��p��jHK�I���Rk��X@�Ih�wMk-��V@�ס���Vn۬�ˮX7��0�R��"H�� r� F�ܛZv��,�K`ᩁ5�ܮԥ�[{w��@��I�{�^ky�aTa�kB�����e]�SY"U��!4gk�b1�
�r��i�+���*�賺N���m��"����Ɓ�9ͬ��f���. 8� sD�p�g,�h��^- �\z���\)])	�
jח�6X�қ�:R	9�A��7���sİ!����4ӆ�%��`�ö3�]2S8.���W�ڴ�8���͛��c4��=/x�6�&��Pm�Q�w`�"��+m��M`�v\oW��	��q���@�we�ځ	��@�L!���[��%$�kN�b��6Y��v1ōq�N���\a�e5ìIM��@"�d@�ben��uک	Hݩ�%z����I�3H��X@���`"I�]����n��srYՕ����	aK\'6�*:�f�x���w�<N^4��α��X#Fڠ),T�%4I�D��&�e�Љ�S5�"�C\�DH����m�BK����i�sVi�F��ӷ��;JH��3��!�����JJ6�$���&�:�DL�Ƿsc��n���1 �m˒��0��swN�i�La^�Mb|L�k�[)�W�߉t	��l��f[�4�n�fL(hڤkvar��D�̖JXd��g�I&[��i�لy���h;ْI�&��;��V�"f֘��am��iT�:� ��c8�(��NH�M��da)��2�&�b��;����j�#�P޲i;�+��F�9�#�&��h9K&�).ek������=�A`M���k��J�QRH�պ͋�"�% �!M���5����@ ����T`�{���)nFWzܛ9Iƕx�Y6q7w4�P�YDH���{m@��0�%f��Y���!�����p��Jam	�u�F�m��$��w"Q�$�L����v�h+h�%
���ہ)�s��UP/3�݉I듂ͩ��f5�f��˦9I��.�e��f�GZ�3�Ё��e������:(�K{��b�,�
l'liՀM4Õ6���(��+�R6Z�Y�@�0FB�ŵ�4E��N�헒�;wy�H�/��V�t٢�Յ��hU@�����wYX�H�x�3�:���=��8h�$�l�ӚKW]-	LYm���N��"I������2�b�11���j'K���]\���Fn�9�MXB�wqČ3�!Xmk%�b�`,��P0VF M��:l�T֖*Q��W�Y��њJL��E����LIlS3���X[FQr����9BVJX&�n(�9m�E�3nZ�Bq�`Mq�H�j�U9��z��,�`W5+�&�]�4�J���ŧTX�9�݇���]�yM�kSmk*Զ��U��_
���7������+{��\�"zn��+��4��ò:e�%P�����*�[cAC�v�؄����0�"�mdp��E�[eh�s�l1́X&��g6\�Շed	�F͗a���������8�-� X��݌�9�kݹa�Kl-d�k�kWvD�;m�i.�!�nۻ���훴7w���R$��k�,p��W��7�Q�7ά8�6�(V��X�4�f���E��;P��A�K(
��Xܬ�bSr��J�ݺM.�:�ǈ�]�m#�H�q6�&�0��ғu�� D"g7��m��[e��mDX"��yHQ�c�j�'`B����z�TJuL�2�kl������ B�Lml��e�HM]�,�i&���ދ�D�[R  ׎%n�&ua0�kz,8�J5��l`*�դ�2:@�h���i*�;v���7{���s�p�D� ����YA9xҜ5�a�8�o\�kZYl��8��!�t*�6+5�w
�BV7h�,3Yvl4� KJ͛�)Ҫk�Df�5�6�2!r�4�ę�a�u���İ��[��!	ǜ	��GwmЫ�� �ŭ��ݴ'��Yݺ����ZV&�՗��S8���-iiem������N:�q��wk�b�7���1"J*�D���h��YH[k�qm�%A�$G.�i"�R ��4+����"D�t�Ǎ+�"6��a��Q�c�d `@�r�ۤ*se"�'Z��&��HǄ�j�u,�N��\CL�Y��Q c k, a�@�t�]o]�/YazE��l����q���]� �k/�����5�%�����0#E�\H
���ue
���JCv������1PS��B1q�"]dI�i��ݻ�"Y���) �)�i���fQ婂0�U��f��t�0.q6X`	�4b`#�d5�β�en���P��&�"���� �1�YGVj�H�JH�H��^��ID�����
�3��"q8�A�)�T������F�^��v3���A��.@7[��(���2��\6�5����	���d����))L���[��#�c
ȬH���L!b�=F؊Ļ����'@!���$��Rgj�j�M�2͌���� �3pȐA�)0;Z��!9�9�W�3	�-��A\	�޷M�R�Ƕ'��t��	�x�ֻf�&�k� Ƞ	֮@�%�K
3G	 �!H���Jx�@�T"�p�M�R!!�#"�ɪJs�MX�����ܵ����y�a	��,im�x[vh1�� emNc$���A�F���$%u���\�v�%��Չ.�����h�	��h�YJ(%���g6K�A��L#�BJXXq4�2�86�c+h�#,�KB&[�u�FuB-n���%2�l�:� }�Y;u��p� �<�i'�B�P"`�L���]�r�̩hBV��h�"j�!#7wvP V$b�]��5�SN)h�&�%�!�S
����!�T13�.�Mi���B:��a�e�z����	���lЫ�i6���Q#V��v���� B4����v쉳p�wG�a�m�K����I��V=^#��*��X�2 m��Mt�l���*���Y���0�3J�la(�2R�K `Z�TDUuB	�N����Bo0��
 �^��c����8�p�b���8�$I˂��Tr�0 mۤ�Xk)U�,H����I�CUR�v�$���:�o3�u� ������`���Mr۶�Җ*4�VJ�m뛆�D�ܦB�u��D��X�KG���ٴ�eT���dE1F6�v�����N%�fo2^^�܀!���2P����5�6�[�H``M$	)
�;9�]%��s��] 0�Ks�{H�Y4�����F�4�qL5� b=P�X�v.�b�\�D�b���t�y����d �4�U!��M� 0���u�#eP��Yä�Țse�ݽ����:���ӥ�� C�labj饑s�!`���\������d���i"Ye׷�NYw
���n�c�&#H��1�Q��l^�f�F�e�:K7�xV޻)nR�,�\*:İY��&��&��	Vl�[�:�$�́G��R�a��%F8����0����9H�%\�)(U�0<��s�v�t��2i���e0�큔��l�!%��̤��D�h]B]۴�w0c]8���m+�HJ��B]��Vq4o�a)�!�AJ��-!ͅ�#z��
Eyn"D�-��\���&��N�a f��ȓa�/T�eVІ Q)j/mٍ�@�8ٻ�(� D��]�5�7\�j��!g��V�[e`DC�g;]4�wrT�5�ٸÔ�9�Cb�,�2�]�RGu:�b�@��K.���-�\J������a���Bu��YSFm{q��B6ؙj]Lm(� �qB�H��$i֝��H�8���:�H��#ۤ�&�BSp1%YĮؘ���Dۦ�M�m���4�&_fI$�lk���.�3`������n�B@�|PT
� \�TX�*H��T�� t;��ߟ�������/ˉ�0���+�}�?������{U�(����hk����X~C�������6g��q����vz����y��k���P��`)�|�_��+��_e��(�4�q~���.~��TK�H?xiLj���_n@��/מ�/��P[jи�>��+4��b��:Y���b۴rS�}�?///-� �ǡX�q�AE�������y"�7��E{���W�z?����ˀ�t�d�YG
�(7�����x�����){��%��`���L�D�	�S�,r�55 ��������]�m�a��}�T��'"����@ӣ&:#�\KeNp:���7f�8�f�I�z���mo9Ҁ�� ��&{��t�"��W���(�2����w( "J�oO��]�Œ5Y�k�
)��J��"2�iC
�i���
�a��>�cL�)1�`:�o2��z���x卡��aj�*�D�&�<,X�<p?C��&)������<�����\����P��ɥW�_z�]��@�T�
��2$F�*��h��1�E��"t�R��:��q���.f�����dj�!���+����r˯:]�f��r�k�d)QA/R�vb�D�ױ�c�d�2��Ovn)���i���X8���ш/P�e�KwѣKK�R3Si0�E)HH�UWLW���v�9k�He��r���x�u�]J����_QE�v^����4��2L���Hېa�<(�K��@���v`\���A>T��|X��!�I1�'!	�O�������!���lM�^�r�a܄�=rx�Żn�s�F��n0na��u�]"�6�%�2��7D��L�m�ѧ�������Яx�X�4Q�i�%�����s�w[��a����̭I���(�֏K�7�M\���<����a�S}��N��t��A�ބWb�6/����5�bLĬT� (�%��6���!���O���̫���'V��MV��M6�\�֊�;���e� �f6�ʹ��
�P�*I�pB��jFHyD�,]g;E�S+�B<٭���Dp�-ޥX!�cM�%Ӄ�%W�$�b�-n��'�ڊ��D,����هb}��0U^�-���X5hGΨ��U�� [�*��p��P�`�I�x&�n�Z���?�u9�6��t�U�"@qs�0���l�S(Ο����!u����m�U�1j��C�8��c��Ś|�%����n�c��A�&��*�t}h��J�Y�9��C�����ӧ��ˊ���WM�$��KMj���e�R��8����C�D�+PB��'����4lh�;Z-)���m��f�y���e*F><kd@O��-݌�m�]��W��0EE=�E�0-1��A ��* �D
�H�
V(	Q��t����?�����������S?��|߿����_g�a}��k��/l_����"�(�_�������1��yAc�G�Ч�+�������~��Rh����9��#!���ȕ��a�~�%����4$�n�������v����0�;S���Y����ؖ��"�S�T����s_�U�W�\���f'��*,�ِF���������<�x�U�Rgni��Rj�üg �4S@�n1-�WQ�u�R��*�C;�+����_&�t�|V$\PQW�q��yܰ��C�Xl�k$	�Je^=f��z�4�8�fZ��dJ�hil�I&2̃�
�t �N,��鞞�����֥���Y��L�"����pªA�D�W�j��� i"�����(�r�½A�����K4 �[���#��}Y��[K�ӐZT�F�X�&���~�0+)��o����(�L���IQ�Qy��I+�i�:�p��N�����T���H)Icy���&����vckɆ��b*�9U2���BJ��+�+ U�������ܦaF��KÔ�H����"�4�R�tur���U�q�J��O{3�l\c���3p������	��qY�m���E�S��J0�spHO�#���i	�/F�ƾ�
 �0Ft�Li/ )AXk@��0��xr�W�>)!���i���v?D	O�E/�1i�����HGE\�7J",=�;cX�W4���;�#�8s�x{��47*j�7��$��(O�׻9;D9��V5=��yO�CZ.А���a>,w�Eu�;۞�1�;���rO�x���L4�#���$��PZ�|�Ɲ��be��c��(Q�"�z��0(��ᘑ˒�l�
j����m�s��[uITfAu��º;�a�����k�w!U�^zhrߩr���V��e7~̀78@�(	��<���yf_A#q��Ǩ�*�/.���;+'���Γ�Ғ���C�l�4Kk�	�e�nG�J�h!{m�p��&��v����yw1#Rv-|mɪc���0�L({\A0.*�:�y	,@���'�t����,���g�^ߟcڭs}�n�kJM<�\ f�ο#��U��:,L�d��>�2�;zI�3��QH��q"�gV�(�+��V�Β� �ΜJH��x�,jG�%jQ�)���4��j���(���Iq����`L����J7hq;�-�3H�|���w���S�$'j0$x�$��[prcSd)dܚg[1c'>[�v�fV�8c�	�:R�#�	`L`Zȧ"0l&���.(g�"0+z��:Yc,!�8�AC�k���
#�L.�`�W$u������]�c����(��  ?3�M	�O�RYq`̿&�$7i03�D��L@�T�%��y�/{ݥ��Kٱ�:�T)�ȖI�|�]Ñ=6��IԎ�RX��d���,[�K�ji$I� �Pb��(QLDܬ���1�4^3��{�#i�o<O	�j���x�t�|[8h*�< �EE**�B��H�N� �Q*
�"" +"�H�HTj
�H�����O��v[���G�iTS*���f) !�j(�F0%mm�W�j�ֶ��p���PP� �N�����L�b��Fo�hޥ�^@�"�T%��ʖGH,��F�`�n(2��UP/2�,��9��M��!����V��uUků��mm�ڽ,p-?ȿ,�i�VC�A0���itCt��t�:kV��(����:m��x���TaL�piK#�P`��`d�U
tKp-�߆T	$+M��l��D0���MGJ�DH	p�%@�0����-���0Q�%�IQj5 (�TR�o�N[��>;ƶ�&��T��$"�I�1p�-]ZH �h����V�T��P&��L�i�ƁpQ��(����)�H��"�$�c�(�)K�� MV(\DҊ"Du@��#|W��V*�m 4� dUC�k��1B��r�ʴ���j�]8�P6�z JAB�jH)��j�b+Al戨`�0EM҂�w*�i�O�EE���u�X�
�3��:wH ��������E�n;���scj֏SX�-U���m��J�����m�nzlmr�X�mE$f� ��@�
Z�$FA�+r�m�_ە����RX�wm����mZ6�TE�kmk���k��kɣՏ'�mZ���i��[V��ݴh��F��U�Z�b�1Vy�5�i*��y嵵x6�����kU�k|y��׋m��ED�%ADI2�V�E�T"�bmW�F׷���-��*��VdLU��`H*� aJ"Kc�;Z�^7�t�ֹV��^-ʙ{mw��-j�,�Se��U�m�mE��F�$�
�"*X��-BR�)�D� ��@B�F]s"��(A*�%�dQ-UjYPBR(�U�E	A@4P( o�E$	@��#"
"�UIb�E�������k*�l��(�Nʇ��a&*�-�ɓ�`�vr�D�X�LG׏tNO0<��+!8޷�c�͝�q�P@������t���# �Ț�齶���x����16.i�qf�"HV�$��%�-@RDZ�( @YT���_ A�D�Q@$TTB蠂�A� *�EAT�AQ�TB��1B�i�&�����O:�-�����f$�,j���Ђ_6gBR$I۷�X�I��]�d�sa�7{�#�]���bf���i��`�}���3��i�N���x��t��"�X51�����]���ɻ�)K
^��'�[T�R�ݴ���
�R��k)4V`n�M=�Ϊ_z��C�ҙbq`K��������l�p��b�G��H.5��͹=�魁��G$<m��,���۾�!v6Vm}�N6�y���J������d�H��chL+KdL!`	8�Fgn�Vq*8G�������k�Xc���cUP��@�i��p<0}�=: ��۬X@	 !�Z�l�|cRsHv�����=vl�p��LDa	V����! �!�1�"A�s.�3T�y���H�g����s&�ZB���{h\�o��x��=c�^�sw�^g\�D�!v˼�gۖ,9�<����=��(n�����
p��'�6J 0&�]�݄}e���lgVi�&�/n�i7Qb���c%�]��X������%��m����t,�@���]F	�$��:��{e����C�Yu<.�2���&�om1Z{]V�eW]ؓI� 1z��<��"q�xy�MY�n��j]l�� (2�i��ܞ]4�����Ar;�=�4�R��B�r�o�`_�H��1�S�:�0�v��F0�ck�47��u.��J��FK��@�B�ա!�q'��{��z��b/_n޲�PWIWV�c	��n����xY$�]�tmˢ�.&���.���!-�VK���7ӎ�e1�����0�����4HB������;gY�VCk�Ǽ��b��!���t)��j�$!�o[�{�� >��3^-&�����q�RC��I@DVG��؛���������@XCR�SH[ۦ� 5��d.���;z픚bmx���/�Й� �cVW۾ֽ�Y�m��CX���u&���ԲmŉT���M�B�O	U�"��
�\j�+q)��i�S"KcrD��9����GP�m�����\ $<�
�P��&��-�:ɡڐ݂���m�-"��q7�f�r�޺{�4�45޲�V`�-km�Hͬ��@��ZJN�X�*keu���MR�z���]�ɳ�.�T���v鉲�,�/�H���pl�(�*i1�dM4�27�&��3��# [X&��<i��(��`�]�]�6��X���,��W��mL��Bi��m�U|"��؂mL�`�"`C����z�cǈ�0��+�����Mw�5�&))L��؅v�[B ����&��=�e@0�S�gj�'��7 j���m�hj"y���N֖��� m�-�$�e$��}�n��YBXDՠ�N^w]&����x�℧���w����J�Y�,���VSL��6�K^�bFS��hnl2�0�I,EՀX�h��|3��N4*ʻZa\Q��ĉ�[3��$,x�(�Rs��/��ԬLHÔ�{|M�'Aie��&��9����D�==d���a�Λ�)��J%��O0�[�F�s��I`{mHCe��ZJ�$d30����p��r 1����-s���b��u�9�D�F�זz���<[�ݼ�B
�bJ+�p0$��[hD��lo�,�[	Pdb��=��X	JXB�m�q�uڪ��5��4	�p/�7Z;�;�Zu�e/����r�k ɢd; +	����� Nx�|�f�&�	��$k���)�S2Rd�&�@�Q���4hڹ��F�4sx�/����Zw^L^Ǌ5[�V�Z�oK�cF�s=v��UJ�jDB��9XR��0�]/��Z��.� �IU*h���+��-_%zV������D�&57��P��r렢���@@
T$$�tF���F��uƉD�JťH2�I_Sz��ʶ�5m�9˦氓t�����l�7wn&(�i)����.�B�Y�Dgv�H9ӛ��D�����.h��$'7g8�ܒ)E�Ӥ�$��. 5 t�"e����z_���a	�������n��z/��t~�͞kA]�~��0uI����t���xt�i����[k���O�})GX�~�F��;C�\�u��-��B��M���ȵ����hH�*WP������C��#r�Ѩ��ض�ֹ�Us�՚�be	����ii�֓6�I �j�ıkU�j䔓-�ڴ[Tm�kV5�mkU�m��Iy����>��H�����]��#CF�P�(fl��PȐ_.���ç��z�U)�4դ�MT��f�Ҵʤ��m���U�W��]o���U�n��6���'f�?��j�E�ת^�^7�u$`��|9�ͻR�1	`�k4@=]��:�ALâU�TRF@��1U��.�堢��\,Q��r��2KƮ�Tb	"�Ƒ"M	a$�1A���e�2"Ș�/uS��bت����m�-���m�x�ū�W3�nA�3��qE�x�ASӡ��'���:1G�s)$�wz��wv�Ax��D��捹b4Z���U�
��Wǽ�J(�㮗��+�(C��ޛ�0!L"���!	d�R1))(I� k'��-`$B��_"�zr+�z[���6K���%`,P���x�&F��э,1��.�;��ϴ�_��g��?���}�_��}���$G}1ѷ���1�K�U�wީ���[�}V>������_V���������e��@a��m���������w�2���"�	KE���Rp!hhشc�s!z�ģ�sL�znb��r�,k�rl�v !IF��Pd_g�}������)Q��5�����M��a����O7�ɵ����woU�����j��>������ݹ�B/&��/�4�WM����kD��g�C�L;
�4�	��_J�x8�;$WK�E;����`?�Ȑ������j�}��k�׍j�E����w��6�"?܍���.]���Mwh&^ut��"1HlzrK$�T�\��F�浊5jV�����\�9n2("D�mrM��A4�ɕ�JH��5%��\Ƿ
��1�y�ʉ�� �t�/-����Q�Y�K�-`O�2��Z#L��Rcj��6���po�oN�Pl>n��Ւe���pI�R�"��g^W�.>q]�_�dlya���l�h�Vd��Tm���Kr���a�]���̺�ϼɽFW*�FjI8�-#��5�����r6+	M
���m�؛��얝H�*PA�W�a���D����qt����ox�ؼ�()��K,D�NP&�gÜHu#�1%��Z����+��i�>S��w����C����_2&�*{��yD6ͷ��RO�}�������p���H�:"�?��$�%�#�`��b9=s�sM?�g���{۶��'��.�8Ɂ��K8�u�_w^�)�,�Btf�*�����Ĺ�Dڭm)"b��'n��`��Ч.�&���h}���s.�ok�*@.7U�f]�s�vR���φG;�:�������a��l�ix�BO�"���H۰ɰ�rY������NCKL�)(k@a	���޲��vh���W��(柆��P#�5D
��A��N��ӫ�/i��"(�)�U��w�Ffd).���H���)8�wƯ�b���K���Y���	Ê�ɻzft�ǖw�rb����i䝍4��ÿ���t��{������:D̸^�|5v���)T9�:~!�3��$�n��T�ʻ/Y.�$H�+���x�n^/��`�O\�־����m�e�)E�[6@��ɧ�J�����J�����u`>d�m����$#)]H�(��6�)��C�y�GE��8p�zl��gx�FS[�
�N��C��x�Ǉ;f��[�ݰ�2e�\�!�#N��1 ͒��<�+�<�U��@�>��C��XORogu��2cz
T��.�-2�N��t�a)�CP�3e�W�K�	�s��9	���o��4�:3<p�� ab��pnE�S�q����/�kd���Y�/>��_��Lt���<���zH�:H7P�v��y��oU���r>M
_�V�@[��-2�.1ox�]u�,~xھ��a� ȟ���4?�^�.���}�;㜷�KLs�B��\�a-�T�"�Gh�g�W'�^MT�CޟR)c�c��p�v|�CP��͜�_zf�PAh�%M��z��(����rM��N�Ѹ�c\�s�˿�+P"��h�9@/(��Y� �-v�዇M�˥��oM�V���.�d�mr��v��R��N�(�h�1ʈ����F�$�̢|���9��e�=|c���;����!�}�;���%o�h��;D�ٚ4]z��?�D�* � �lj-E�nZҫ�T�B�#2I0T�2�^�D�$Y$a"Ȇ"�	
��ITh��k���H����]��"�P�B�-]�#&��d��f�ͺF�� ���4׋�
$�^wY6�zm��Eo�mr65X��-W���׿^,�{�H�.��O]� R�Ȋ~�ۤ����bX�﫟l���Qm%�mE�m��S�n��%D�rj(h��%�x�9�E;�QQ��䁮Ʈj#�Ճ�U��h-�+U�[�碽��2E$�1�b=u���0���yڮZM�[Eh�X�Z���U��e 23z��<qsrdҊ��y��;��������>_{� B� ��k?��?l?��Po���o��?S�-�_b�{ �a�Pk���{���B��a�R�98d�A���$l�4�� ��g$5���eH:�߾���ͱ׬�i��贬c�#�����m�q�L7����?v�pX� "MD�'����u��7<E<&����@|�S�T��EZh�Qr�j��6%�c�?�h#����܀қ����!_����V��,�,�,ް���=IN9f$�b"
P_D�4�Gt\�<��0�ԶB.�p�A�[	����A%V]"�xG&�a��1�rT�=����T��N׌I�2��$wa� ��d�<��Q�,�ѣ,@ �=2��Bcp��
��+.{nz��~��뮹r��$&ps�Z�G��?��eÂ�b�|<�ꇻ�M��K��L��B�V�8��f��;�p���ȴ"9�0�����,�c5j,Ȣ(�{-�Z��^</O���K9��t�2f��(,���t��ZD@r�o�#r���$���p��XD�Ɖ5;Uƴ���
 �H����AW�*vX��)��� ��j�ɥ,�$�lQ�56�a`�H��3�3�N8��R��a~Ht���e+!�H��AB�e�B�R% �k��ҷ��*�i�#!��u�m���1`Ǐ-Z
X*N\���Ƙ�e�Ia�%8�W�NS�g�kBY�a͉ -�a]�:hZ�9�'�()z�7��x8�Ѽ�i��j�22��-TP�-[,T�4�GW8�2�<i��a�xU��{�&>?������*3�}x���a��|G3��/gC�CAİIC�x�����Lxi��G�=-2DÏin9��Q��19:[��!m�,-����.�1�S&�Bn�:	��J����$)�U�Un�����ʮ��X�� T ^A��
ȡ��ͫo�kn[V��E�m_MW����So;�3j@�H�Fa�<�sFƍ&�����ko��y�ӥɔ��^.A�6J4��Z�EoW6�EQE$hԚڛκ�w]��/1�����;�H�B��o���6��V5� K�t@��	F�s[�Dk��5!6)-Q�گm[��������wr4��s��A��MslZ,UclRyܗ8�;p�wE�K��b�I�\Ԛ/nED��h��Ph�*�cd�������[|�1)�Ƥ�JlA��*-��+�Q�j(�-��h�<nVJ�ڹb��LX ڒ�TT[�rɣb�ƨ�x�F���\�nm��뼱lmk�\�o��-�Sk�*�U���1�v/��*
���Uv�_
ܾ����ܻ�ߎ�֕��j�QUF-ŭ޽]_�z]�F��5�wd�9s���b��S�p��j�t�ۛ;���]wiݮ��nm2�Ƌ���)�]���э�gܭ���q��-�]JtI�@���+%! bĨ�����1���6梺nwv.[��]ܑ.�IS������Ʒ.N�;�B�Ycl�� $p`*@�Ǝ�����'w���<�\�wuswur\����$�6$�n���Ү���vܱ�:�RF@�$S	��H��e2DlrA䳺9;�H����k��]9��nW9���|��B�AE����*��IR��+������?���y/9��C _����������z��É��X�5$[�o~B���$� Ʋ�I~���?���!9g��������>?c��\?�vZ�-����,=�����`�>o���?���~a�O�����Ỻ�k�ms?�Q�����'kx��_���W/�l2�c�a&��!�չ_+ �'r�T���v��$��P摑#!�`�T���K�S�� � ���#y�M�S�,U�R!�eZ�!kn�=����߼���m���=}���n���R�/K� B�ZQX9lY5�Z���'6��+r�Ek^,s[���k�v����e\��y!��b�\U����~�d+��b�+ƴQ�Q�W���^e�4Uh��uz���kۚ���m��u�jLjƊ��^�6����m����ոV�(�Ɋf4X�E��V�kW�o�E�-sەX�,Z5�-���hئlh*.UsZ5Z���.%%E2J�6�V-Qm�Z���豲��dٕ�Q��zmmr�đ��TV*)-�[���ᵵ̓H�K	��]&W���FѶ+b��5o�o[�skq4�d��^��$mF*K�mcmo[἖
G��4�X��IQ�ܺm\�zj-x؋�Z��km�i��ƙ�l�i6(�(�m�j��կh�媼�͔����P���W�^+�o�x*�6ە^ըګ�=�jXX�%i�/M�,lb�J1�j�^����{^�(�nE$�&���ӝ
s�E�Q�Ƅ�ms\��֨�U�Tkn�V����X��IQ�ـ�ъd�65ͷ-�zZ�V�����q�Q^ܱͺd���M26�&ƍm��b׎h��kh֣[r�i��7��Q���H��4N��PU�F�ѭ5cj��j�W)(��ʞyy�<WM�n�D&�%�&(�Q�h��k���DBEN� &()tAX!�#bѱ�(�|�]ݫ�J&^6�С,��r"X�[��EZ6-��ŵ�-�6�Z�U�nh�K�#$Ԛ1�h��1���4��BƂ6��5�o*��j-� �˸���� $�L���#!�F3H��ƶ�Elj��V�Z�^���j9��&�+���u�,���zq���6�*H����A�T��_���ڽ��	���rƂ�E�]̢�2#d<�ל�(��:��H�H�Q@���6�kr���V�L,hۜ�$\�W�1%˒Q��IdB ��R�W�]�I���cj5F-��h�+k^�]�y��lmF��l{n�cS'.�4E��;�hFCӢB��b6fCF4C����W-kڪ�5�-���լ-�Xѵ5x�H�5s@Q�cX"�$̤�)��7wRE$�×�+!lj���mmcZkM�˕�oJ�^�Ƣ��K&��71˻��d�%
%�],��n	���%��3F��zp��}?׋��������������1�Q�VD��H�]-
����Q3��C_OL��]בZ�t�WYm�m��&yk�S��#m�$�6�ٔ1�5˨��n�.Lf(��t�n뫼���{�K�����_��ݼߦ�w�}�e�9N��<���}���G
�읝xOkaU>ER$�ߝeK��}����/�~.k��a���e�����K�m6fLZ�B��E_]���5���H�Vo����3q���1�o�N��1q���{�e?����N`�A>�?��1������g�z��]�\S��3#�������H?C%�Y	>VXQ]��lBS�^ �#�_j��Sy�J�,>�������t��#������ԧ���%o�؂�C�V*]�}̙�񨸚N@ḹ�F��Ě�c$sJ�6����7�H����}'���o�*���v���A�T���15�c&����u�`���)�ȠSdcJR�E|��|�]����[���������8u��@<<�6�4��K��_�ԗ�#~��*��_��aA�я�7Շ�Yø���G�ԃ����/���/��}/|/>Ț�ߩ�~��\���,�9�]ȁ*�`�l~!o�����}~{h,F�fy�����������"9ȡN{���<����@��ĕ�T��O��ċO�^~��)�_#,�B{���b�%8���H�6?���3�ñj�J\��'g�GP�v{7��<L����"�F>���s	wb����?6��{l(,2��T�Jtw^0a�x����}$��p�sW_+Z7f���������1e<\�so�ԝ�AgP�V�1�qz�ɟ*��r�T�]����)�Ϫ�v3Xlҷ�i��v3�5AE�g�]�t	?	s�#&��%��G����3�d�</��>tN}k�+��w5��	&6����Y����;���v�~|��<�9c��֭��~b^L޳�P������	9�X�G7!1+������S��|\�A�"�C�)U$����cl�Y"<A�&�75�	_k/{e�$Ì9#�Z\�Q�t�z��|����
D?U��U{��[�ﵖ)&�S4,]�?�O�q\�ȋX���|��n�W��MR�ks=��d�rႮ��Z<� �{Q�/�#���}��~W�F����Yr����+ˡ�RMl���,�8�m�zut��+�tl[{���2w�[�u|�
!l�R��G�/J�\�� �GKt��n���T���ʘ���u=��(�<a>�9#�$��2�_{S]�E�1[q.��xF��?-�4�tյ�-��9א�k�M�&^		.���k�lY�x'�$ (lY��K��O9WL:ҝ�������H�
�_v�RJk gʜg�CoE�ų�Ԣ��Ni��׸E��FVEd+���#嶞|TAo�9�M+�/k�9lSwb�*wcm�Myaŝ�(��w��ك{�hO���:�Y�9�15�mu��	�A�Bq��n?b~���D���~��a�y�Dq-����[��[����p|�io`[�!�W�"�#�� ���/ev(K� �t�����.z�+�I�_	5�w���o�q���A1k�RL���Gs[vT��/����AP:z���3������C�*�����l��Zq�tNTݸHu�}⋗�?�6�r���q�-�Y�v#�'~�;��5�p�+�������f/[9���o/md5zx����KN(Zs꿇St18�Ivc҄b��)~6�/:jū���f^G�ӏo؜k�����6�S�W]��=F]n��JOZ�_��LՙC������`8=\�Nz��&���x��C{�z�PP������Y2m"Tn�� �l}��99��;UƳ�T�H�ڏ�e5|���� �%�p<��@ <��6~ߎ�;�m�����N���Z������nٺ]�s߽�>�J_�{�N��O�;����1�q��������������<ףR���i?�R�y��ĺ|�n���h}>��֌��?m�~��p��u�7�on����S���`�����]^�ʿ��P����d7�GH��� ?	ʁ�ɝ��<�3�I��?�*k�x�=!Y��o���}t�v�q��l���-�����I\�m�� �pC���+��m��s�0�ښeĳ�W��� �j�[��R�ǖ0x S��L@t�0��e�j*�)K$<�X�	p�e=��T�?���k��nx�vǗڙ�9i���|�eGz׎ʼ�<�ƴ�zͅ9D
�F�8_��[y� 9��:��i��U���� oa�=�͜�%&Z�
�2��3�8W��0e����ap�!���$�\D�0,L�'ʷ�
W��8K��ۗ�$���Dl��I y����jQ��k� ���A�,��~�G�8�F�g~,6nqӭ�`���W'8�nW�./T�7g�j#-5�v
�5!3bI1C�����ԡВ�	`�4��4Ч4�HFt`�:g>���o��a�ǺE^}��u�I�jB͵�	�3Fe�Չs(�`6#%A�Ll`p���-��-��-+�
-0Јt1�Q(8�B���A=�����=3�AE�J�$ElӃ��A�PdF0��	r�X`��t�\�\5�ӓ�	��p����%�I+�D �W���M>���5��)�?xkT�:Owg� p�7k����8�[���p�m��M£9pi�RjMD4���,�W+��Rh��p�v�78���<�y���\ţ�\B$�8cR[Ů�775�F��Ey۴h�).m���r���b4G<^$�Iյ�Z�ݯkb�%%I�)��@Ȳ B �Hp�������I$������
 ;�� �Ɇp� ������:�(!g�c)J��B��W)�!	VM�*����]�D���b����]�PT�"r��22�����vW;N�r���\Q2E��
BA�)'9�;oA�&���	�}����coA����~o=�OM�=5(��$���OK/�EqI)M4���Aõ�T��TT��-E�5��ض�5����Vت�Z�Q* PB���d�R*� �#b� @`�L��9_I�W������g�l��?��$>��7�}���E��w��?�z���-��I����C8������>��Օߕ�g�/��G�*�?���Vj�NOdk��+_Rٿ�T���X @�����	L}B=��� �Z�:�/ Y�ʚH�{�[��o��<��=:>c'����h�����f�t���sM/�\D�Z�1��C`�]z��6�   yyy  yxT�hǷ9�5hu��Y�4u]Q*(y;ߵ��ig����;�YntU�Y
#}eq�8�c�*�,�-�y���!�xDaWb"�����A�K��xv����V淭�>�9�"P�,��:�\��CF�DRg))z�ѱ���-Wڅ��m�bk+��]�[\R��S�:m���"�����R�}�Z.!RӚ�����e����,�j���E�,rv��! �I�#+�8X#�.;��&�&J�E��dvQb�F���t�����lփ��T1���˥:T]���M�T���d=s����A
���8�K�v�9X�����	ljp.�8!�I���]�Lꕑ����d��+<�@W�+�� �4 n�U(��y��E��5u����[������HA�i���)�	'�6�
'
���S�U���ts���l����4�������"t���w�C��yR��l�zUP��*jw'B���`�$Gm\r��:z����>�e�6ϱנ���ٳ�;�����L2l����O��&Yb^���}�-V��2aO�,t!�^2��Z�Df����oL�x����ŜV��8��F�Z!�o�.�Eh02Rx�Oe߼�ڞ�.|�gƖ���C�Xl�'��6����f1�y�7�I�-���ǭ���v��|{��e�q
�3��jkP��^����g��^9*�kFC�����=9���fu�V�َ���R�2;�b���w
V[�i������Y0�� �˸B�VA�7L��*����k����ش���=2�)�+�7�F2�1� 9Yq��WA�{&Z�7��/QΜ�.�s�Ѕ�ue �s�s�݂�{���p�S�î��3U��9uf�CohX��πھާ�&ﾌ��b`�#���^�mi*�2Ak�GN���P��^E�E����ƣ�߮�lbqۃ�pUeo����A��Qy6���k�+R�l�	�V^�H��6�' �w��00�#����>�i^}QQ�!��B�(��-��AJ�����_ù�v��

�����2�9��Y�Ñ��$r�AD]�*�w�Ek�5��veD��\[����۫���	9H6�.$��k��r^cnU>ْv0�H-�V&��EKfo�(z4�P>j�蜻��А�$���
Ȭ�9�"����9�`�|v��D�ڪ�ِ�Wˢ�6f�&���N���g�
zb@˱g��&*�j#U��@�:,!M>*c���|��JU���+_���5v��8�r�j"2 � �;�w�7����i�~�8�y���cﾗߝ/O���?�R���������4z���>����p1���V�����}�Q�?~��6��e��7�_��i�55��z>��O�xt����{�;��?���8��^�W�Z�o����z�o�@��U[j�.[�?;e�eH0�y�N��7�!w������
�rQ�d��	N�!�J�2L�ƆZ�=���v�1	�!C�H�ֺ�
 �.��'Ŭ��Nw��Җ��R^�L���<!��Q��G$��*���%�1*D�8���8h���h�A�=#�Ҟ~|C�C��ژp��׹�Q%��fޅ�$��"'�m_��J��@<�m� L
:]�AgeÇ	֊Ր�Y�,U^S�� 0�+
\'�l�2�M@lG�%sŀZ��!nPX��l��A��xr,Bb���q ���Z��C��Q�Fnbۂ��Y�b��ؤ��8��0�[�@�bR�X�L���dA0��q�*��������<y�A*d6�wZ+�`3�&��:D+�v%��$�9�Υ,�L�\D�Ybe>RA�f��"q��-��P�|A�V��C�wg"�s1�6�� �A4��C�+�3��XND
E(36q͒�Ь3)�(�S���X��J�Q¢� ���Pg�!^�|7a��1���/_�-	�����҇��Q�3���9��)�	��1�E&��R�Q����,,	��09sY��m�E�f�P3�P�ؒ�B!I���aſ0�DAP�T)�[衛oR��l�ǔ�
�d�D�H$Ă��Hm�Pkw����mn������o6�g;3EQ�"�vs�-��U
�?oe��U��~��z�!�2��W��w����uZ���2�'�Bv
�l�BA"�@C$Q�A� @�" DX����8�����txާ�á�}W�u�>��tWp_U}(`�?+�|�[�������'����i��vW�!"����3�ܷ�J�y��Ayyy��6�![l�&�b��I�O����'P;���VK�N�����~�b5�@��������	)`��{�n�C!�G��w��q��̼����8����� ���[��[1��;�kX���!l�����Rj[1�/���d/	��<�.�'��a���t��[6wϏ�9eM�ݯR�!�)����;ѓҞ����%Y������_��<wai�ܯ�����Gk)�"K\��/;���p�� ��f�MY�[-��-��i�m3Ԝ�<i4��!\��g��Cm�-e����(��P��)�0�)��a��u�R���]�cAM���ϥC�-�A�����6M�v���h&�a����.v�^s_�:J��S֒�s�^�$�-�Ԧ�]�n���C�s���E�$�x��%�3;��خ'�](�]�U��{r/]��z��}����8�,����L�]QH�f�ӧ1-����_~��b3����S������K�@�[2;f����/;�X�dW�Q��
nNX�P��=��\IX��%נ|a�"�耷<R��_����f?'D�uEWXV����=�^֣�ehMĤLDd��?D�HG����족��Wm$��픓����`���/-�ͨ��B!���Gz��\�
v4�.o�h�ڈ�dnWq:�&�pҕ�X�'�ЙV*��}P^���NC�'A�ߏ��uq�9��5�Gdqzr�e��k)�@)��N!�<�I1�{���_�	�����fƻ�|Ų����R<g�X��z�C�
�5�翯*ɮ��8B��r�~�s���gK8�ף��<�:8�����+@Yݷn������o���2��x��bT�­���ً�F�u��J�WC�lcJ��^,jrE���g>u|�#�0�D ��woc���)�b%{x2��f8���Ap�#Hj�I��44��.ь]&���S�pL�h/*�x$*I��Gr�D��B�b�O(�G�c���`���7�/A4�-����c�5�È�\t�����1�6*�\�|0Ӈ�O����$K���BO�G����z������_:����Ke8�X2�lKyԛ��Q�C(
{K�&�<�������Y,���z�烼 �S1p�ϗݕ<j@{�*�S���D��]��GqD�w�~��E}�%8�tH�A¹e�xT0���JqCD�(�FX��>=���8:-��~|P�������>u�ejD��\e��9\�K�MwPЦ�/�_͌�߇����i���9�Xy�[���C���CK��"�-Y��m��Vś�uEeP�׃��5��qO�#�u����P�w�q��ⶻ�oY��Ύ���8^��7��E")"V$U u���麞w���O���6p�B��_�s�=n�����o)�h�^�5B?;�gܼ2�4g����'��M(@���� k]�u���ΑĽ��+]�Pπv}���:�bui�iu�?ϲD2��
.�_=�hZQk�3�2�.� Ua"�]�鐓%2���XoR�0��%F+����~p��C,WQ���@*�$�$��-hҴ@Y
�<�g)�ڙ��(�>� ��Z�)��fJ��|o�/+�\�5�-ϖ񮼪_ht_Ǖ�׷�-SfV�5�$^1ۜ��hN��������w������@�>������"��K6\ ùI������ �x�Z-g��+p$����XCR�,��%�i� ��]T)��T�V{�VDA�PN�p@�0�8@�K��f�ۿo�me:q�ƚâ��玊�v(iu�k�G,�R<�C0t�T�F������L��I���g�6؄P?PI4�Dpa��+�X-��y�%GX�K�Z�l�uݍ���iI�1���S���M14��&�s�!�(�	:C��ŗSUT=�2�H�0��K!P�(�1R83Ǒy �GD�^=��Q��6���Q������:K�_�<�!�L~�����ڤ�OasT �@�I �d Yb�)f�� <0��H����
��� �UE�p�d͵�oRR+�I|�=��L��n��9c2
�����[[�� ���rKFF�M��4]r��\�h�61%�����O������?P��(D���p�w7��������5�=fw���=���|_�_�������t����S���	�y��~��=!=RF=[�$a�/�/ �z�������5g��=+"+�d*�����D���>�m��2�Q�-ҟ���h�]?3�E��z�yظ��z�G�ªV��,���Β$[���߅)�g�33Id���L��L;��>�C�+}n�@���?4�i�A|��]˳?i��n�4TQ,Zl�/��:wf�:�o�����t�ّ�-�3�<�o�������y��:�k�΂D	�z�杂Fn��Y����˵U���$�	Ps}�G��������שz$f��m����^�1'�I�͸C���֖p�3C�Sx���\�<��}Y�q�K���:9�u:� ��%K�Lvw�qy2����,�Z��=ļ�O߂��@�ص�]�uƪ����Ií�8WGe,��w��W���%<�/����'I��:�HS��).�$&V�^�IV@%oa}�$�4e"H8㝥ӧM��m�c��q� �����qR<�|Ʌ$���[C�?����]�o�]+�x�M�$�p��mq��hOF %;�G6�2R�|݄F7Q�ҝY�6+N��׿��kG �-�NA�p�����|C��;>ٲ��.�3#Z;t�����"OC�w�O�?�[u��:��e��-[�`���8"+U�>1�zi�a����(�u����`�|`B�*U䉢�[˜�a3���g,C��0;>~Yx�6c�bb��N����5������Qa�g��&�.]���9ͱ$x�8]�����V2��\&,َ8n0�՛�`՗�\�[=�u����A�&y�憏q�q�ߍi��;�K��u�\zI�k<|/T8v����������y��:�N�C�Ee1�U3��⬸�Ď0'�7Z�\�n�����)=*H�4�IA_1b�{�l6C�K�$Jn'u�p8wV��X��WY���xޞm�ŞJŊk��ˋ�HR
d��JAz�|�4�4
�J/�T�{^%����؍����IחN��>�?N���J��� �f������N�4��L�m�cm1H���{]i=i�@u��,Ud9P]�S�&���x<:�,�7�BϮ�V��$R�Sa"Bֱ�3�Q��^e�*�L��o���!E�5����̍����N�;|F7���scj
�>�	�ؠ��
�(�m�74a���b�1]pl��3a�m�nks&�	�d��oF M����!R#kp����xk�E�x����G��[L��|A�ߚ��م����s�7���GsG����?4]z¾k0u�Sc �����5�1t�C^50��?5�ӧ{%������&&R(9��-�aG�Lh�-
�Ǯ�[Nj�sN�T���<�!�����j�Z�;R��/�}#�>�'���d*�MD~�)P�޷�jQ I��y�2���t��V �V�´*s�F�h�wۦ��,mM��s,:��R�t�G�C��@� :�#������ϵ�{�D���B����6�@�H����9O���D+�f}�a��� ��O"G�F����}����؆�~����}jf����������w�$s�S��������f�����;~�����-�e�=3~�̪7_�XK7����'�X�]v�}+�<}~`�o���q,��4df"�E$��MAN��ʬi� 
9�K��V�J.D�e��3:,@�ek%�S�i"�(Aka�$�]�;����y{>aݸȋ���q����Ц�������,��0P8���98�:)���&ߞh��@2P��140FC �k�R�L���+�BHjM4������H&��_ ��I+x6a�� �Rh��;9#H�|s�=sH���ఐ�&ޜ�}y�g�ǐ�g�N;i�OW��r}��Vv��wp��m��uy��Ȳ�9�y��G}��K�n]��{w[���±����R��>���6������|kF��Ӯ��7����T�� ���l7�-�묃�E�)8qݮ�R�MH�BEbv�:o�S����>�;�r:W�\r�1���9�w����}k^��_��i-�������O-m��r��2���8�I&ӏk��K��
R�p:*�ĝK]���0�Pj�H���$$ VZ� 1i��1���mI���[_m����?s���d��R#ռ�_.s�����~��������>�U��7��^���=�=�n
���U���՜)������Sx&n&/?-��轉�A94Rq�6�*%9=�E�]��/+��wYWR�q�k/6��0V�Pj0gUH�S	���:��ݸ5K��sCa��Y1i�=�*��0���f�ڥ5]6&iҺɊ���A������1]�ڲ��̡�V��av����w].���@Əd�lۈ��,��}W�b�{�cT�v(^և�<�>e�[����<s"�'�n#oܗ����c��7p6A4adgN���V���P��X��}~�y4��b*zu��졢Բ�CY�r�:�8U�oxk(�6�+���Tl�B����S��bۢ���˻�k��٭ث��{��9�K�#����V�d�U���p��9�����;�nOn��X&"�Wu`���񬝩�s/��A�1W��Rs�r�FX�6�x�O�i��*оgc~?o�+� ��s=W���y�K��.���[_l�|/!��je�3��#��>G��F�����KЇ���Q3L�C��s��_Z/kꈁ~�N��=�_ �����1ܺu_���� �z6�aЈ���0��1{��$�Y��lz�\�ٹ'�Y�g���P_���3�2���rN���G>׬�(N~<�R��#7`��Ak�d��$b��M7
�Wy+>�@ <����|&z�D��tu..3�-�1�%jvٍ.0�v&U�<������4|���Ӄ3LG	��~Y�w|O��Dcx3.�d�^���0����Q�>�S�9�S�.����}#r*�_�L��N���a��Ҍ�U��k��o��\��%|Ё^\��r�E�����f�=r�i�,q>��|�:��iX/^1w�`��8�m(R���!���<UQȢ�w�Ã�6���1Z�̄tF�?+;�|�{�H1���IW��XqYZHq�{�1�77t��N�l�2�d��j��9�w�ŋ�_*@�G=+���S摘(���Ͷ�+�<����=B|mgP� ӑ8x��cl��=-��$�#�h��>�c>AS�v��Cu�/![��J2`��K-�2J���2�6�2��N��t[�D�v锂9�}`�	����*p���Mܡ��ԋ�FĨa!�=�X��������et�H8'yU�"l_��m������o��q��q��u�����;��f�Z6(���>���9'F�.��U[��N|㛘Y�i��)�OM�7�~��q�*��6 �M7�s��<F��@ڈ�]68{��q8=�9^ZLOx�6�&�/-�bD�P?�;��ʵQ^Ha46�������cnuE�׭�����/9�K�q*��=�N�Y]�G�7�(���L�এ�2�D���`�NсJ��#S7ɓE#����W��6@�\�Wm��m�Y���{�Ę��ݩi��[��8N>lM�bL��=U6S	��`�2;��*���V��m�<-"~d"3���4���@�����l��t8�����Z�Fv�ϟ<Gܽ�����;�.h���wJ\�*��r���eQ���%����Ǉ)!�1�����������MA��EL��o>(��p��Z�ӆcOR�t5G�� �u��p`,��CNK�ܚz1|�<v��Xc�i�9���	��p�d[�=;p��H�\	���T}���]Mp!82Kn6h��zV5\(��E$�c���i�<d8���1ju���p�a�1.[�´��M5H�K[�ͧ���WwE,��a��ˠ��˶� oOr6����}Q��I�;�!/�N�u��d^[u�>�����I��p<�E��^4�YK�~��V��:���*|��p4�T>����
D��8�4mC��4WB�=����sN�J���mvpkϠS��zH��f׎Q�߼4��;�i���]Q�����T_k�NvM��e��G��}6��t�N�M�ioW�:��d�]7�Ǖ���=?K���s}E�kl���O��_��;�:���~�����;��i�7�����<�o�	����'Z�W��N�n+����2���0�{�}��zp�_o�x{i�ø������ev�f&5v��>���-x�{���㣵���������{y{��>�S��ƃ��~�zi������C���,�o)�����GAW[�9�nuX��O���q��6�pw��W�]�3y�t�?�>�o�����>x��߮x;���/_�w�]��1،���q����xT����
�;�24�B A�DP�(��9��x��Dቂ^�]�z8܊7��L�"�8
k��#�����U�����P�}��9�bF���k������i����;�2�;��ӿ�n6�ۮ��V�|��u�$#�ᗎ�:��"�/v��s����K{�덼��{ˍ,�$����3DH�,�"��� �'5�4��s�{$$r.�.����=�>�;x����v��?y�Zw[A��=h/�>?o;�Z4/!�\�Hz�=��^�ǧ��oW��ӷ�|��Hkp�i�Z�^�֬9o΅;(QYtZݪ�ԜѺ�v��Z�i3��z��F�[�DZ�5E`�6�޽'�*(�+�?���OY���Y�;\��9�y�S����=\���������d!)7�b�	}&��1p��	��90�;��]FD��^*{@�O=�9��Ұ��
�w�L��W�8�+��U�d�ي#5�����|�=t\
����q*�M'�R���<��
��o�c�����W�� ��\�Z�wGz�v�7�q��!KWL�[PT�a��/vD�\��v�Ο&Nq��F��@��3*U���rn*3#T�vH3خ���^1P�[|�)�O.�\��;Φ%�&TC�SYu�5B�:�Ӊ��{�]�{G*`\Z���Q��9�"vb�&�t� �U��
�@{��յ;!�ڗu#�l�a�/ �u8�Ό�7�r�x���{�n'�oo/'r�l���*�,Z��o� ���#r�a�N:��u�(�[����}�6#�Ov���j�B�}���93"���i3�;�m�ٵQ�f��vȻ̓�W��f�������|��]$��bg*�dƷ�yV�ׅl�뫒F�#��Sэɠ)��T�ռ5"�c{�-����ߴRt*� �ǘ��ꏵۦ��=�d<�5��!-��v/�w*�AU]�`s��s6�U�d���[h��jQ��Y�sw�:=F]��{t����.�O]OLv���O�><�����r�W?�_��>&�����nW����K�s	��_�]��2�5|�E��7�J���{��7��N|y#X�X�W���ϋ����[�N��J� y ?Fߕ�>�K!���_��[eߓ�������4��-�_$��1�c�O/��8dO�3��Q	�՛�ۇ'�Vם���H9��O����u���6�*!*�c����;6�<�I�5^T��/���Nܾ���j�����N���P��l1����؝q����Y+���KZ�.�]�_���u#�-ڔ���h����9�}8@+X�%��q	��B|7B��*^�x
"��Kv�Qsn%h�q��T�>/{��y���㝊�5��Z�-�y���hJo+�����&xk��`]�c�'��)��b��.}����@d��p�27z�W9Vэʤre03@�$�ƝDժ4��o@�f�!^r�ߢ�,I&��;�ScQ�����N1��=��d
܍��JT�0����G��N@cˏc([WR�I��Ì^U���Ox�����P?u�k띶�]��1C�ψ�L�T���^�'98��8�QG(B����ޒ��󴂱^�XUXA4��T��̓�6�i��-�{gu���韯�jQOMA��pt��gH��m=[:&G�a�x��L�jX7����*-'�Cwm8��v�4
̿�Ⱦ�7*ng<S�D��j�E5d�܊*v�L�Kre�i�����#K�v���}%ɳ��40�o
�כ;_:�'4�A�r2n;��d`�uX����X3@�d��9�gv^P�$�N0�C���9b��!�q���3Et��1�d�eL����=o�X���t�W~$:�v�Z	\�A�<��"2�gU�E�Z5q�Sh��\C�D�=+�,C��p2�Qf�Ӵ���ęx:&l-��CBV�s��-ws
�����,�Q�Fc�-4�G95G��@�'����tw��r6�ׯ�@��J)*U�:wK8�3�U�����J�B<aWE��3%�7�#�ei�0�3rt�1汇fÆRU_1�&�qD�&��!�v�������GK;f�}N�f���"�(�ɵ�ǔ$_QS������}�E-čòy8��U�z0��2#/ay^L�2I|y�L��ڱ�d��|0����q��i��������HĔ@߂���.�}I��B�(��㒻OK�0��Q��$��_.v�\��=dl�ߖެ探��?�Vݯú����(]�J�vq��3s<��T�*������pd�Q,�b��3�GE��{�!+���qt�!�Wp��J���ƪ�C�;ߪ-.o;�]�U4�y�1�M�{qv�y�ft儺��;�,�=G���&¤��Kjݱ�l����@ �w
z��Ea�}&�ʷ�S�T�S	��*������s�aN=X���^[�!�]�0��C%��pSW�-�����4@���C�4{�{Y/7I�ZG�=#fK�LX����֩<N�wZ��~�՘����� ��x_��=E�Q}�~���c�������7�ج��K:�*�>�E�/� �vqm"3ze�X6v�G�G�N�~_���B>�V�y�ǿG(��唉}�J�;��$!)o=t���ˍ����C���u�[s�:�{?�������u篟�����θ�ƞ�8�eVt;y���[.sV���i�a}�4Ɩt���'5�_���\��=~+,ƻ�~���Y�|:͢J����{u�׶�5�6����zl�y��O�E���09la	M8�n�a���h4e4hۄ��|��c��%��׵]��F��o���t��6�w>��HK�=��%';!�s�|�%rp-ut�Pb�o.�:��R�>%�����/������4w���n�_�;o��>�~y��oX�}�X����[�o������9���䰞�>�6���¹�~�RY��Ct�>��u���{ަ�ִ&4d�hQ��|����W������[�l�:w�B M���n0m|BE��Z����T5R��䰑�W��M�m��_��v�g���^���Z���~�k���z8��uQ � ��Q��FV]ё"%�6*4Acb����a<ڠ�$H!X�H,S��:7�������x�G����������_��D�G��}�Ov�� %6"1=E=���D������mg|�B���'�G�lrX��p<����f[��{&���e#1Bf?�MX�^���z�����[RkE3Z����Y�4�� ��>Ы׌iD�f	t�h��"��Sָ�yyyp���@�@ %�a?�a�k	���Q|�{��*���[+[^x7\_\����+>���<��X�
�rW&�ĺ���'j"YL�r�jTZ(2s����.��+[�0b\*�BiTJ���Z �V�3n�n� 2"�TLǐ�m�O嗰I��ݞY�Mc�yz1�S�Ќ��#*z@}����R�Xsk�M�8��B���jUQ�w�x�l��i��C+;�O~�pT��WZ6*�L/7cҍF����z�����	������0��h�H��OV�6⌴�$\b>�d�2�
��Q�-��� ����p	�V	L�v%Y��P�tLff9��4�D��=��b|��ᣧ%�e��kv��'HM]|�T#Uvi���h����4�f�Jo�o�K���d0�-/n��g	k�1~�`���Om�e1�*�p�/��ؙ���Dpfұv�S�'�,!�G%CÜ!(�r!#��)�,���f�vo�FDkeb�8��2F���*f��Ȓ'[p`��"?1��cxQ�~�B�K�>�FU�>p�h4�W��C���<�h� �ڒg5�`�c5˭�VP����jzH�5��8^�]���W=(��t�F�ny9� ���3�m�b�.dK�0�O�_3�TI�6t�@����WH��"�#�����3jH��a��I����5[�:K�}�v�&�縓uU�:��q���⍌�Co$�{��p.�1��h��E��k�Ljt�L�0���QfFۋ�E�D�T�N��+�W2�׵jl�d��«�S@�!��`� �@����n�Y{a&z�ATf�,�(�CG��R���D�굼�#jxfR�s�+g��CK�d5L&n���i�խ*ԌJW]���"���e�2��՝��β�p}�?C+��&N���kX��(���S��M=�J�>��݂%���Ny)�]����[f�Qg�Y�4æ����^e�CHM�mA��\�O�ϯD2�;��d�́8�m�TDۤ�b�F� {��Fι�t�����vE����5
���2�G�ӏH�u�iO�s2uBB���P{�p�S�=s�=Ǽ�(NG��DQq6��t9��^���fga�-@X%:���j��c?d��6b��\bG��"�d��U��\85,��l��Ƅ�_,T�.�Z��lT���6��������cQ��R���pH���c�nN��-`n%A f�(=�
�Q�NyZ @t8(�6�E�?�8�瓢������>��>s�������q
V��=����c{�ŢAX	 @<V����|c���=7G�u='E��3�@���Q��o��1��c��o�5������zg�\���L��<9�+n�+��ƽz�}f���c,/=#g��.m�K�ϗ��}�Ow��ֽ6�s�ӌy�j���!:�M?_�朌g���b���l��]�%�����[l7�_���(�/Mp��A�?����V�Zv��ް��wv�f�.�F��7Hqb3�4���+����%�s��|����x_F�|?=��h��m�z����,!�m�����w��������К���������~�;��:翧O!�o�괚�'���A��gx�������kbw����ҳ=��p�-Gj2��[zR�����/�CK�Üȇ=�Y�x􌷻U����+s���]w���8�XF1����o����֙��d�^�
4����v�c��"�|7m�~!͑|��)�����~�������~� ! ��臠D����h�o
������r���w�G���O����G�4K�(G������Z�3{��a��&*ǯ�c��l��Xi�sxq���u\�T9My�r�N�$dEv�qO#��1�#8�4�T�ɸ*M�eX����n����݌�y
٫Z��c،4��j��Gx�Mf�����ﯹT�C_nI�7�"R����M��#�^D����F�թn'7,j�=6i
e���/�"�qo3k�毱�/�k'�73zr/0t^�T�:��3mSR#a)�3��5�8���<�Q��%#�;ʼ��F��\�wj�i��u9晁��+��J��G>qW�;�xND�����48�W���t�ƴu���ؓ}]��*J���9��dD��[�b�mFZ**�\+s��a��g"�+�.�����)dM���W^��1d֞��w+�&�{��'����*��8o٥��U��\D�r�T�+�q3{1�mL]gnf��k�E�N>v�S���M��$Kȋ��MF�������_ �P�E)��MT򗽫�gU�L"&6���㳻��otȱ�&��9�.�:&�+fj��X)�{��iU\a�u�im���A�R�\�[3�Q
g����R.��ӛk���ۙ�1'�6(���Ė@���1v�K}��E���v8"7ˮݻ�ov�!n���CP��Θ�X�1ױ�4�z(B�� м�{2UnVD�*�j�.�Jܵ�/s�˭�s3�a*�ʱ�8�j���-�\�҂���w[S1�y[z����=�Fd��H4�;�����H�S�wYQ]=xlȣ��x�`�����k9�Pe#}}t���I���$��s'�Ϫ+���9���Ω�-ќȜ��FI���������\��1}w1bȝ�B�m��]��͚�]�TW�Ӽ�Ud[��(R�/`��YPw�k�3["I�v��J)]�-OY���W5G\S�-���UwǪo8�2U�ۧ�4��>�5��[jc�=��ԟ�y8��/1"/)��Y�,����̴�g��QF�a�.�bN���z6ʻnd*�5Ӡ��i���9�j�GE݊ܙ}
Ǝ������<W�Έx-��/r�l��9�P����.�Š{{��&�K�ET��{���:����ґ�_���
j�r�3�ۏh�/�3�Î+�`��
�:������<箵^����1�o�5���UԹ�o�/h.rE�Aܕ�[�ү�O(��ó) ʉGZItM���En0g�f#�eH2��<�ې��{�����^�60h9�3�n�#v�j9�bO,3��IZq�n��\g�����V�l��t ��j,��.Uc��'_bqkz6D����yVʴ�����뽕�	�}�������ns�Ld{Y8=�s�h�%�T�27�kd�us8�yJ�Q�Ӄn��{���MTĮ}���%�܃Cu�Z�63M)��0+��}�qڊ��D��2�PB���mIW{�PW���w�[1�tg_�w�n]������[�$ˌ��)�)ѱ��˩9�T9)�OΟ&�OoH톦� l�}<��pS3{���(�C"pmdÔ�NP�'-��|�*8�C�b�l��I����2byqܭ��X�0w*�.��VQݽ8S�r�VFm��R9�����"o�{���8�F���|��Z��w�J�3Fj�*k��]��s�%�Kͽ���,�	�u�/���1�Q��Y��\lMS�l��Nj֊�is!�n٧��QԔ�r��pZ�[�y&v�
�Evl#B���Z����-M�\�an�m�C`N�yw����vcv�a��ݤ킂I�F���reY�s4#��t�n����.��gw�^�Бާ�.ɼ�B0V����O;NDU�A���Q���)���=�h���ŵUV䛗�2��8��iz�,�vy�w�v���4AW�U���u�C���k�dlp�C������弆�gNJ�����:�HW10Dcj�<o&,�2b�\�����Xl��l;�[
���%�	No�f�`c�7o�&�^C���p��]
�
��t �}Q�]��8�T��m8�Q�5ĉ��;0��K��;�W���Kʸ��븩�jEa�����ggaU<�0���E�}� ��\�:�F8���50��)��KsQ��=7D!.�Ȧo���D��5H�|��9�'*V\���冶���6�S]�o�v���MNb\1�뽫�q
 u`ʍ�*���47�W@l�A�9r"ʮ��eoR��LQux&�P؝���U������dfp�&���j2�M
;�w��3�L�%�����5q5�:5�cq\
qs�L��,�ܨ�&�51x��K��S��,ӳۊ9m��Ac�dk�їӂ�pv�	mK�˒J� R{�z�p4����q��M<+)����-��"sg2�e\�,N�4��7Ě��@�}8�\�OHa�v�lr�5m�+��5Y��ta�����®�wy5Ckn"�$��轱�3Ӱ����Y��Q*��0GA�����\�˦���~uD9���tt\�_�S�5�-��k�x�륊NB�xgsɻ��L�wFu�d��(@iE��ޞ݂g�m�����l�6�iۋڑ�ʢ��8�OQb��V���TD�a��2��C�ȕ|�4�3�lMk�q1'���ݪ��i��3��XhC�y!]��ڨc���7Ekۭ�N��F1z*�$>X2�(�1d�ᦡ^�޻
Dl�� �bb���o�U~�rS�oo,���p�N�ޥK2}����X���gk��J�r����,�s�3}���v�x�'׉N{�S'c,a��)�/$6�R7f,���.1���B1�v�5Z/�˴�P���SHd�4h�35\����׃_����MV�ul��'G�2�Q��a��}RӜ�Ωl����#;�^mɈM�'wn�B[<LeWu�E�mI���X�v���9]9�&E\r��X6v7�^����꼷u�[��U�7;�$�loX��lB�|�HT�x4��M�J闆u��{��ʻ��������ڥ�!n���s9�o�mW��
�A�q�7����MA�p��m���vpF+L�b�ȑ\��A�&��Z���&Z)�K���'gh*�=�<�2�u=�F��;����Z��F;��vM�<4��ЎX�����af��t�v�I����*�����z�v��T)ҍ�VByGQ��aL��s{$��EYvw28Eʪ�z�\,q�6+l'<��1s��*og�֦�z/�fw]DK+a1�aw������<�ka���khwK��ͅ��fS�/��lN�͹��סsٹ�}�8��
y5gff&B�'�|��Έ9�z�õ}N����@��"nk�7S;>:�f�U���w���Ԛ�.�]�����{yt��n�CP2�rBs�%YQ�.z�g�d��]���*�eމ��ވ2���\}'�S��2�Q{�d+��UZ�x�vM5qy	R�î.��7��v���gU7�Q�x�"��x-�,��	���Rȇ�tNu��^������OD_��u���
,��Si��<9oMќ��}R������u�_z��Q��t��A����7�FB"�FJ�麮���V[�o6�0��%|���UL���˭N�>�^N��R����c�ll%�r$�(uq8x�q��F�%�5=�Ɂ�7�oǪ�輻�Hs����び5(r�����viθ�!�2��q�=�����^�W9�����4$�������[��s-񫬭��鉓�$вr�j�޼��էj�=R[��s1)d�it��i�nnq�5Y�ΈP-Ø�1ӽ��h�%<To��b�zwuW��Su�[��v�Me����K(FzPQ�}�r'�:�Q���|�5Ʋ������r� Ћ7�]�/N�>��0�ۈ��ҪzN�D��}D:�p��c
n{4��Q�j��p�ֳͺ˘=T��^X�y$�m��W^8�I���o���P&�k�P�n�[�2v�LG����7�ʚ�˒��APr��qG�Od.�����Ot����}���'^*���#0�4��}Z,���Ģ"���v��$��s �b���s�E�wƻ��ڧ�H���ɚ].�K�'\�
�Dl`nY엩ʎ���N�ߒ�9��k�5�N��UQ��� ��q*f��'��ѕծ�[�
k'
�̐�z6�f���;q�L�+b� ��Sv7�ki��Ȏ6�c��.�gN�5O�AΞ�1Y��0�n�{"���	RS/ޯ=���n�W���cOb�m<r\&ny�Js�*�>�;�[�PlK�R&gj����q,+ܕ�f)��*�E��[��._m'7��Q4�nmk�1�fq=�Ce���`��"�cQ^�ہ�뻵��	lB2&��gD�Ύ�z,�OFXI�N2E�a�Y&�@գ�Ҡ���W��K�W��h�*�5��<�<uD��rTp�C�-�9����K�0��G^���N�d\�5���J��xV����N�+��plv$���'B��<�}Jm�9V�FJ��Q;�*�:���pY����Mؘ̄��6���ߢ�#F_�C��D��&��U�s���7s���T�5�}yê.<�}6goc��7uxg��^R��hR�u�ص���
���
E���˚�YS�W���ޕ�V��$��MV*[�a
���
n�/j�h�U,O%UKsn�"�uG:F�y<��󺼬���y�[nL]�;ph[t�5r:�,�����2��b5�,�VEѻq�t��|'zl��J:�Ӆх^op]UJCDDH�7WG<fc�7o�O
ڬ�[5�1b��9K�Wp*y�+��H)�<!Ef�93/�U��gN���t�K���y�#��ۓ�K�����5d��pr5vy�Y����^���|���D�yϲ+�5�5�w1]��=�Z���f�,3ul�OGos#3Z��:,�nZ��s�X�6�:�²݌1淦��LD����s��B��]X��FK�d��<-Gk�v�S�㦰j��'�n��T�V%q��o-y)�cݻ�d�9�{4/������"�qR�]V�1=�������y�:��K#o"�ٝ$��*bm#��؛U5�c��uj�����ۢ�MDٹWt��[�,b*�c��r;�=D���2μ�6+�㛋f�*&so*�D�d�K�pe�]�t��WJ�uuR��{bi���/!au{|\L��3Μ�1V�Z�SUn�}3Q>�V9�����;��dE�v�T׵QЪ��h��qkk+�5����L��m��ķۉT��=5s��>�ÄDTt�9������9}Rӵ�J�̗*���2��ry-uө�2�R�yS�"��W�;&#��eŬlҌ�ʨ닙kD5�|�}���NLFQ`�6+p�D�Lm-�5d�܃y�[EwnՎ�����Yu��^_	�R��AQ�v��4�x�(rj^��ȮgyY�S�x$G2��=��ء����f���h��ʣ�"a+����Klog��f����0�[��{�����t���ż�'C��u�8wtɲ�j�w����;��2'-U�ފ2v�i���`���.�u��:I���M��ң,�A��5Jo�̊W#�������7]��r��]*�gL"�r�N泮w�_^
k�o������:���t/�mU%�v�MgHXP�"'��sq�t�j˾�1U+w,Ֆ��w^ԓ��}�W8��l|m��wquuQ{�3��,Ѷ���t7ɫ�Q6���w�j��Kb����f�5�W=-�{��f��4�K�A�UGa��S�oj��!�+��+����&E�6���4��f�F�F;]��ۮ�����ȳ�Y�G*�R�⨽�="��N�bY�\�����7�i>�f�ѩ<7�+���Uf�Z�`��9ٗ���z+��ٕ6)N�����hte�=�U���T�8�S��v�]E���nbJ��֢/#F��F�C아I��z�Ѷ����]3	��s��޷�tI��ӌ��RYv{j=r^�I��F
ғ"צ�m�wu�O!U�4[K/l]�:�F�z�Y��� ��D�*E���G+�S����\���v%����V�]�'|@�׷$��$��s}3�%�q������"k�ΩS<Vte���l18+��)0cʹ�\���+3�ξ������uv�KD.؁��E���L�=u#�{�� ͩ�*����n'�j���Ξ��VH��r��K6�D��˚J�x���w'9VO�Wf�خX�Tt	��:٭�s��N�{v�6H�]��(s����ޜ��4f�s�ڻ�c����/��D�CB�S7UlV�=�*z�m��ow���j��T�ȊB���'_E
���3����i�LIӱ!�co,��Z������l�:�i��9:U��3�;o��2�љ�w��h;
e<ܧ̙�������ȧ��0E�ݏh�Gn^�R%��4�|G-75[�ĕ�+67������1xV�6��������{���	�眳�m�ؼ�����ɏA�O��[�l��q���u�˾B��*���.P����*��PI+-lK���aL�.n1�۵��r�*�%Ä�z9*X3 \ON�y�=S�Ը˒�
Jr4,�H��u����^U-b�^�kk�l�����.]c]���;��1��qw��3��NWP��b�s���.�k�����=j���ܚ��n���v*:��ͺ9s��GJ�1�+L�-<ܲ
�4�2y�by�Sq<�!�:.��k��9�<^�r���P�:}1�eZP}�5���ٹ��F�Hvo_ZSTVL�ٜ3�wOO]MD���4��\Pe���H)˫��3���=��bQ�iLJ�n%��4��JU1�6�M����P"�'�4:&�(	��Dh������TI�H÷�r��sjϮ2�U���75f��}����%��o=-�7U����TgN�IEL���;̙��C5ڼ�=HV��.�"p��2d�-D�_;w�ŷ�wF76��b��q�wD.�9�`���*#��͙�v��I�WaQ�{�sy+WFG7v��<���xw1�f^�ӻ���9Vcuv5gN��<+��<\0f#�r�8:�魉�8d)�;�"�U7(�7�+T�Sۿ&(^�c�]�r��YN3�c\̣R�-M�J��[�Vp�h��l�u��Ƚꞧج�ќ	��afș��9pTgo�C��@���F�J�w�y5�e�E�4̖�=۬�sG��Oi���U��D�_K涖�Z���ʉ�* vuu�j*$ffJ�=j"V���w'��屭�m)p.�>��ᛰL�ܝǧ��	�Vǰ;��-%�&f��M`K�s$��*�,ƣ��]�9��uxEE�c\wTFLi��K\*�PXOz��*����������U����6f�fp˨�F^�7�"��r+(+�N�����[6�1a�8wz�*�4�uvF�4���L4���w�}t�5��D�!>��UsP2�E��+#�aPɊ�R��]ے�,�-e�fϽOV�u�&)U�vl;+or��ڭ��L��8T�[��}�u�c�R��v���_�fr�N{b_�n�ǹy&I�7�'�pa��Y�dLWV��;w�.�&��Ns��na�v)d�i*ڃ=E��Y^�jm7\g��љ����mL�xg�fI>>�ͣ����׼:o�b/*n_{W�����ڙ���7%-Z:��ԌC+_^���@�	B�b��9���q'��^�
h4���j��ͫR��e?o
���3}Njn.9�lE�����!��ܺyUX��.��uo��r��蜝�$��:��+^f�p+i�[r�&�v��w[� �m@�'�������o`qix璚[+�n*�X�_Y���V��OZ�����3�j��<{�V�nY���&bou���y����`i�J tS�u���m÷�B��4����Ѽ��ϽR.vN㡸6 =P�k��G=P�]Rp��̻Ǿ;�N����t��u]�55�O�:!���*�.�l���2�n�J�q�P���&":{�.!��M�n7<2�Y�q��:�Yo���>{|-�!%T��<u�Pb}���U����0���S}$�ʡ�w�$�KoS����({��=��Yo���~�#C�s�;������\T�k�Q�f�e��D��t�ʝ]'sܐ��9�v�&��ݗROyѸ��4E>�ф��ז�LF��{1�Z�j��9��9�m�����.zAꚈ�!>B�P��q��Ѝ��[tL3����DJ�����).��x��J�5O{E��Y������XP)nf=��8o��ʤ�����&�f'��.�K�����X�ˊ�����x�S�n�A4v�Y1%�4�̹�uU\f�U���W%e��Ő.j�G*���6t��9��h*:��'yP���v�Ed�T2�Q�t�ڲ����E��_�_��k�sZ�h�mR1�kC+IZY��v�.��Iœ������WM�t����(��6����-(���3Y��2��vfѤQ�Re�1E 1��1T�"��$,�IEM�����c��ƹ�n�&4b)#wk�I!#�d�2iLn���7vwWf�Q���&@Br�n��76�s�	K��:��.]7@�f���u�Y�\2F\⢹��]q����۝�i���X1����7n��\ �.�4��w.�I(��w\�w$�&����'u�#FɈ��s#��ݎ�!���7K�.\ܮ�n]�w]�۲0]�hwn[�M�qbKb�-p�F�-s���ҭs���� yyyyy��������˿�y��^�����~���Ǻ��z~���/O�/��:j��O����I��b|f�`O{��O��O��~�]��(��|4��╰�
}2��R�����{�x���l=3,���ν�8��K�/��/K�E�|��E���۷_�駋Ϛ'�	ȣ��o���f8�I���/V����)�#�iP���W[��n�^@����#�+E�+��o�H�����^�xf���h34���B]>zÛ�W��jH��I�)Y��<<�b�D�֍�&�N��<�jUR`��@.�{�Ϣsl-fS=��J��s�y�=�`�*_�"n�ZN��V�ge �9q�����l�H��78I#'��K� ��v�d�.$�7�����i���o��f�����|ܛ������ے��5 ��:c�*+FQh� y�3���n������/l`�H���F~��-��&f]U
�i�v�)��/��F�i�˫�u��'U��H�b���?�����
y�go�r�14^���5�#�"����{r���n��3������ �L�kr�U{ m�ۚ�9-/o�^6�i>w���ʨ�[�Dr�I���H�G#�T6�aғ��C�r��"\!�\���65��0D�ܰ��^�a�L��Vu�4�Wg�\Q��G�;{��x�ơF��������S��J��m��2{třѫlzΕ�7�4lӨ]5���e�)�FJ	2h�����좽L@�U6/ZHw�5P�\��^�Cw�X���T�PE�b�M�Ǵ>Xx�zUԳ�y@�7���ٓ"�Վ�pܠ��F&���=���$p�S�Ĩ�]��%qj�'X����\<Ö� �9��(I��Ik�>vɪ��B�/U~6������μ��9�Щ#�}�lӘ�)��s���Z7��$y5l���'?����'1�VM%�+�X ��
1!�u*�d�]�p� 8=�fi���w7{^��F5��9�ߌ�Q��=�518�:^�Г�	ݜ��q�Y�!�`쇁��bx��g��#�vݦWOCW�p.�h�u�F:�띏nw�L6�6����%�>�Ą�
*R�dDwp�YP�L�P�-sz'A"���·-�(���t�4�Cƣ�*W����	8���«X#�'IA'�u�����y	~k�p�(�2X�W����{���u��惇�B��A��g�0L"�M�eth��3J�Wi��>����Z�A����ֈ9�J�Lox),���1���*���r���Wd����$����A�g��/B�xRNh�E<��I�����%�Y�3',K��cʡ����裧E�	�D���~��$��%a݌6�t�x�;�,w�FV���
f�.�۬�~''���F�nS�0fa�߻}c�)'��A.؄��]��Pt��A�gBR1(��Ю��ʙ����u��f�'�9+�y _�z�c���|_f߲��5��n�������?��Am/I����Wم�и� �?z�LG��
�X����y�{:\b�[Z�[ZS����6�!�U=4��u��<u�4ߏ%{��M�4��'oM�)���G��tҲ������s��)5������ć���������;q�v�^��xUӾ�����������h��zw~��m.�rݵ6n�9�3m�=g��*�0g�9�X-��WFt�Ƙ"�"�p�e|�|ܻ�c���o'mn����48횿i�GXֳ�k�����h��9tw����.���q:�gR��ш�Ut��W	-� �I�}q+ϤUѝn�x��{�n��۞�A�%q�>JFXtȡ�Q�hI(�=��j��4ڮ���<�����v�g���w�8����D\�
� 
��x���=߄��?�s�C�s�VgA�<?'���kM�v��g3��[��~������ܯrg�e�D�D)���|r97���2;������O��|S�� ��s^�H,�*�cBl-"F�L�/x| rώZ���-�ii2�F*�S8��g�5�����2���5�Y��V�pK���܆bmu���$m~s\f��������-݌l#�p�'���  �`��~>��C	t��������2��3`+�7��}�E�FFktˑdj�}Q'K�P�#d:�4ކ�LR/N������q��3�F�9��Y�P����!]e㠩Pp�:5Tγ�2 �4!ej.�.�Ã��tD"�Q���e�Ak9�I���P��4-��^���|���!-A�kjԕj&6�Ҧy�� ���,npED=�3�)/�6���8FW�Sg�N��1�I��G��翆K��9�nW��f�||{�^y��h��$��j�"�&�u�UTS���_O���-UmǷ>�)F����P�āӜtW�*�2ބ"z�o���("���<��{�E.�-�n��_C�iQ��U�K(�����d%�tSO�gċ�C���cg>��J��=$��Y�rW�M=����_Y
P�g�3�𧚛��At�V�$9�ܙ����͛�b����&�5�]W1S�c�#8׀���I�^%�/"���kw��!R�~�3�%���1�S,aD�C����YE�C
�.��!.����9Q�@�cfO���ȁ�QS��g>�s�e3�-�d�D��^���[��f�M��ns:s�A�b0�d�J��ˉ%�-�V���Ɖ7oK�ZrY!�"���b����uz�z�i�M��R���9�v��n��n���.�j�M��P'�aٝ���g����'d�"*��-Řy��
��'M&2^!5V�^*`[�E}w�����5��7��v@իc\|&�u5g9��'�2υ�ʓ�uH��8�֭4k*����JZ����"��^I��f�ҳ�L�.b9��&�/%����l��˦���)U�欥|�]�jcu|�H~pV32��X��Y�������><M�s�x�c�#&�;����*_/�"iR�]'r9�6�R�P�D�sZ��Xm��o�4�)�e���*�n���S���t��Px/n0;�B[�WMj-GDдk���@Pâ���X�4S�^�����c^��6����ռw��R����zn%���o�AQ���ӽ�N�����5d�4pb��"z�|�w@��au@ac^^�ρy0�o�+�P�OeހHbDҒ�A7s�y*N��]�"�V���N�J���1\)�a������������a�uy��>�C$|�l$u�܈�uӏ�'q+k�Ñݢ�Z�9]	�-2�u��Zw&k�S�n�<�rc@�WuH3$8>��$?�B)�$GF��Sa��>��ciJ��hk+Wv�4M�Y� �� @�� %/0�����K�C/���Y��,��3��h����y���6�ۊ���8C�\���S�������U�%{�4Z?�	ᆮvqn],�ʙ�1^M���#��G:��*t�a���zmn�C&0�'Y���Ѥ��AYb�s�gb*���A}�W���9���ˡk}uۦc�Kc��듯@�C�β3x�Kmy��V�Mq)�����������,.�u�V}�1ݞ�>��D���˴ڜ����[.��h�͖2i�D��\a�*�^����/ͬ�Ơ�^]TA��s+�3��QѤ�I��u=oO�����C��s_��|���R�tP5�����Mh�M}]1B��FR����m6���.�c�ɺ��c޷|���i�1���j4�O6�j����&�2p��0�h���H�S����/�ϛ���� �+n�}}����'���4'M�t4�ּn�*��]yZA�h:��=�Xi��U�ewZ��W��m9P��2��U�f3�	��k-��֥у�Q��eR�@�C��G����==:6+�ꯌ�Ī���}*>��j>Z��"76sƢ��Y���U��<��zn����$������ok������i�}߬ݸ/���&���@)"+P��Rʷ���jʥi�5Ml�-�VZ��KiZ�ʹ����ݺ}[�eI>�b��R_O�%H>�>ӝ���T{���.1k,�b��E1FS`4��"V���Z����8F-���Uޟ~��%QQ��XÕ!��5��W�M��cz)i<W{��:�4�,Y��&��Ø��b�s[ghY�=�U�i��a�y���$�� z�@��7���y!RDT�X�s��Nf�����zݧ5��pE@� �b��H�B Aʊ=�u>��Du0�+��6�AʩP�R�	=ĹK8)��X@��5ue��b��nuU�q�J��G$�V�Ld�����|�4�'��PU�h����%�]��PQi?�0@/L�Ѭ,�@D!�ŗ_#o��6��o�{�o��w��|��������jZ �P
" 5�|����D��yxz�2�*��;���v�_7��vv�4!7h�Y�i�3�ՙ�a�t�'��YgofI2|d���؝/r�W� M���9�}Nr]�"���gԘ�a7!���ƒ�ƃ4�� �:ݐP�����bJT�UDt�#��J�&�)\�h%`lPT�1:�M2Mv hR�J�n�]ck	���8��E(�6�O�$���*Bo|�$� 6����4Q@Qmax���5(UQ+:O�X�F���.j�X-7|fDHI�����A<*P�RB
����.P�U����򠔾.�(+�(�#��}H�U ���j�b�B(PPՄ�� D��)s��0�HH�כ��YDP$KB�8ވ���y��+$��#�Փ�J��(7�*M+N��'�o�b'��}��=9�⁒8��	]�+��	�i1)w��P��9��j�G��
���J��!-5��g��G��0����&�/Ơ@ �M�F�|N"�H�iDm���MH7 �l�d�0�HJ�� {�\�H�P5�ڰ�
�:&R��+D�2�>��MK�,�iN�$ �TJs�����P@�EW�&p��RUB#�E����GW"j"1񚜛�܄��0��*Z���)��0�:#Q$B@�	�Q�m�TI�v��҂�R �@��KM6��	�:��ǃ�r�b�$m�e!��i�o�@�f~�Ȍ�(�ze�1(HJH��S�R�n�E,@�	3$���u8)��&�r 	b�B���K:��2R�2}�I	@$vP�oa̸�H@H�Dԉ���J
P�Tܺ��T1
�F=F܈�
@t:0��\�)$rg$�̑���̀(���5k	�#�@h�B�`@w$IáH���=!ʇ@�I�	2	��Wc�ħ,aP����J#�T�F_S��o��de�p@ʦ�)�d��X���j�ĞT9�7� ��QbMŪ��T���I3,�m"&Rbb|;�<0�(���X�F:��2Z8Ƭ,jj�5��)e
*VeS}Y�_�<vP���.<��y�'�v�<?�Ӣ��{�vÂ���?TT0����~Z��: z���ay<��5P����i�C��i��UP�R.U$��/x7`�
��8J �
$dt#K"����,L釱�TYE�ń�b�
�ԣ�rE�T�Tb��2���Q�+Vf1X����(8s� R<s���<���1fk�B�m=A(Hԉ�A�,��Kɻ(b[���5��"
�  �w�v���n53��a�Lg�?Tя�#�n6��@�$	����O���	'��I'x�lỄ� �H����Ukw
}=)>����A��wt�I�`ʤ��Qb��4j��n�v�H%&�f]���R�	�޴S1��{���,��E{/�j@�12���"0��2N� ҡ@1#���P�T�*�GI��T�c&c�or`,�i�����0�/�(�~|��b�!!=aG�`��퐑��H��H���Ǣ,}��c�+��|�g��(�O��ˀ�����,��س*�N��I�	�����'E�:)ϟgt�e$�@t,IL-uS5�Ԫ�2�FD��G��^Gk҉$��65h��>=��!���(�8�	ݭ<X:n��U��5����� ����AdI1f��>Y5fɰ��_3����`�)�!� ��3,�֧�6��8r�L�9����<?SR�A����E�0i=�G�P:!A,�y9��໣ʪ��+4,C ���[D`, "Hd
4">Q\��RA�F9���=�FUT/X쪃��'��Hv�:3��Aic�$B3$ț�؟�ԔD�Cy�C�L��`�I����OXhm������u)6%�*��;�7�_��P���1L�U�)�E&A�ʢA�o�VD�W�i���;F�"�F��l��� }�w�m QD���>)�H@ȷ��%:D���򕹧3��2Vz�+>%z�.!H��)7�qh�f�$h ����6�a�Ȣd9�������c�0[�P�K;!�$|0W��V������ʭ07zYD!��G� N�'��Jݢ��;�� q>��D Z�+A��)�/��
.d΂в�@��qd5QWŖ�N])��X;U���q+Tɵl�X����{8�l3���J0� R׼t��P��X��2i��^TweB�щ���e&/,�eF �QA4���"(���e:���D<U�ʪ��(�-�����(���f"*��U��u�qz
^h����n�k��Oyőj�s�i�ւ��!REJ��C�����I�TD(���a�=��%2�:-�xBZ2��	U7_,��u&.f��˦\t��^K�����6�X�80 ��#�O��UbܲK��V�eP��UBɔ1'�ϵ�I�$�J<޴H
�R��T�H������{�r�+��{H�+�EG��$��������d�*�k��jdj��j���+Dq��� ��Y���� �Rb�+2)B�g�e{P���oڴ��vr
'I�&��0��Q\�r�<1a=x��6��C�&���𖄋$z(fR���,�l0�`Z�!ё
1��w�Pu�����M3��,|"B�/`���T�1�VF*���L���˶���y�2;�$�j�֩)���s�F�*��N'���!��!��V�kdM�	(!������[#��|��1-����>�&���)^�]��t������&gܵ�J쯙�0�3��.TQ~)���1D%M6-���a��\�	��51s)pTc)���KВ���e+�gC�6��qGм%��e�g�1����<������[�^)z��. �ʷ�"UI� q�򏷥�$�ĉc�W��?=�iH�E��ֆr,�.
}1ү��QFZ�j�#�[V�[����us�@r.\��WHH�ҫ@�q1ƚ$��Ԝ�h�;8<M`$ɠ��>��D^J�3>�?{�n>�$
���$KԂ(z�I0LT����qZ8:�q�iZKƱG�r���� P�Z�E}= �D	FȬgh2��E��h͍�jT	V�7�iʤ�V�+�|�٢D<AC�Bn��w��1�@�T�8]�:��dH��)����:�% N'�5���{��_�s�C�ts�j�Z�Eg5B�.paWޮ��/,K�6/��A� Y��e��)��$�`R(l��\3� J��b11)�#����¡.*�ŤN�<	ŉ%ʱ`X�껭�d:^����I^���$�*��BE&��&L���],�����PEC�EC�֝	�l,'U*�d&���JL;���0��Q��ծJL@LT��R�zع�����l����,U&A4eֹ)��(ȉ�#���v��ɨx&���6FS-e�OZ,��r�C�\���4��lUh^�sR�1JH8�"r[���](&@�ɂ	��@J�������|�=k�&�nTI8��3�S���}�,L'���P�bE�j�B�Nb2��h�>s_j5�J�Z99*,F'9DJ`΁���̘<_�.T��4�(f�3R_0W���r�K�vm��n\Uپu�^v�X�Dpe����nڠ\��{U�\I
��-����:N�[(P�-L�7����&�i@K���i4��M����
R	����S2�ԇ+���$���l/�#F���	z�|}�\����B�C>�JBjB�oP�!^�❪3$L�4faZIKne����aX���়akj ��ʖU<L���	&SyX5�����H�e]&�_??I@�J�t��qlT%M
&�s��P�Pu�E~9����đ������xTڏ&HF�e���;(���)���\�^@I�	<�Ib).��ng�Q��BE:�-�x,\�Rbǥ6��(�
5��7��0�����%�gW��&hd����Me�Y$�Q&.��D$�"@T���&��������`)�,ʮ�,'Q��!3&T1p�2^�J5$���3��"��	�`\�0�W��A��B�=K`B�\;��6P�����`���&��HOS@Gi�A*
�	�����nj$$��cY�e �B[4H��+*�4�̢D3��e�X�ܬJ(�����$��٪Q��H"�l�I��u��WN�5�G*�u�|Ҥ֌�^���n�>�z";3�R�KZ8(i�ȗ=���d]hhK��:sx��d� 9Wg�*c_�����pmK���XZ����	M
hk_Q8)��(��PJ*�[j�+����Me��������H�X�C�Uh!Q�p �h2�l-�c�K����P\:M���LN%@� |�_p���7N`iQ�7�ቛ�8��,��ҩTH��0�
�e+R"k��w!��j֮:��^u�Z�!h�O$��X�V(��2���d����Ⱒ%oEd&����Z�S$�&3Yݧ���i1 *)0&*'Vee�|��W�y&�kR$�u���"F�7$�*0&CImĖC67��I�Ϯ���Is`+��bU���ɗ�eBC芛�y�����KL���CE��f��I���`ʋYֳ32�Qj5h5�֪$�:T��/��*�-���MJ��:¼��k+�@5��ƭ�y(Jl����DL�j�P�,j-�\"h�PR�U��b�A�(�'4�0�u����Ԓ	j�'�nc�)1N��*�D�h�&����5�P��U����9����J
 �U�D�kP�A0jA*M�PR�k�#��&Sr�7I&Z୫̄��bQH�i%H�ӊ	�C�!�$۵RCY����u��A�"$��!���v�t�aH&���VSzf��z����.!��~ lk�o�,��P� ��z�/w�aU$�c&H�%�����I���F#�u��Z� Թ���JC�RER� �2cA�@���(�e�����s`� �,@ma�Ð{frp%k*����&MMGW %$J��$+1 �i,�H�(
P<o`2hqVi	
ª�O��?R�P�Ē�m!��$�D��R�{�T�q�[K�ir4��W
�(��;-�ܩ��2��T�5��(&@��	���j�Aa�$ytV.*H�l�24�f�X��B�بЊ%��8�D���� RDT,���Nҙ@��,�7��"z�%h�Ԇ��j ���P��*�T���# �P�q��]�đ"e��Aw9�g��������a��u$��F\�$-@� bV����ab���
�r�n)s��`2�E�"��F<�A>MP���@�<#�DZY�Ȥ%��WQJ�q�6Ć��9�q}ө���T�A(��i�y�DX�r4(�+���(M��3 �)tғJHV��P�&3��RMO��H�H���R�D��(�T�)9�8�4��'riI"�f�(f��.�}V$!{Ô�MEF1P0D)J������x
P��V)HK� Đ��M��ҽ��R�ЀH�b��q�ا��H�&@��	���D	�Q �9�b�Bq q`���E�@�)�D6��	r��� I������\�#,LPF��� D�6�QB.dR$!BV/p3jh�ԠyuT
j℠���$� ,fQ!�Q�U��@&F�Zi �$$
'R�Q8�<�ruaJ9J8��� �fE�PؠiL(��	@H�hɵ��GX��UT.'�")D����B h�����1Օ1�	" ��Ԃ�s3��Ȑ%;��?W���~����k4H��`	��"#b�U%�H��!p'AH�T)x�8��a��E���2T2��0C"�Ę�H��~�tI��+ Is	��i6;MPuY���$�%&���DK�q����$ՠ����^��
m|@��1D�E�!�B�	eR�Y�!�T�L��g�x�a:|1�9���,���6����|U`j\C AN$]�dj�DtUL���9xlM�b���X����rT�#�r!-�Fd��P��B)#r��TTJHr�֠B�>��T$/QU����ӆ|����J���n�YV�]0b��RK���P�[v$�D���H�-T��f"4�P�¬��c���Ɠ �U�j0�Z[=#��br&�ȣ�K��TI�4Ŝa����*1Z���A$@��bP�5Tq6!j�,��FAJ^]#ս�G�W����H���#&fZ�-6��J�RE���`��LzQĊ]`I �D���JeŵkP�Z5���v*h�@RH���/�h�>)��_����풁��*��R⶙h�|i�i��jmR&�}FP�FxO�bB�m��諮"L�������2�F�ĨR��4Ġ�(��,�
�vPÅl0`Q<��Rd��y�i$Հ�V�*�&�B8�Z�I�2̳��F@IC��DTU���Ŀ~b�(l�T��h�"��]��J�Y�K�2��FF���]�Q(+"��u�\i�p�C���ė`R����B�C*��x|]������X>�-��m�Ԋ�*��PN�xd �M������jގ�*�V������j�(��Vb6�)����CA}�}d��P���h�LJ��4	�(�Z]�g�_����l�Ћ�.W,�"7�I��6z7�T���E$�Xo����)`�D+2�n�C�SNn#G>�} �(	�n�x�c��2DGtOǶO����(���#T6+3.���@�|K�(3�����sT|�!x����b(gX�Q�J�[g-�.S��N�X�6P�>ĉ_{� ����E��N4<�ȅF �Y�q�c��b,
T�fNʵxQ�,�p�ǻ���_reUU�Dg��n�A��Z�����$�%�#	e5#B��f�#%��@�������7�PIBނJd����R����1pf�4q\٩:���C���kG�+�G~��?kC�9	��l�˵�^9�x�8���l��+�����JP�+8ə���H�7˭iX����-��b��]�}୨���Z�C%Y�)$u�AB�z�
b��ؗ�(WF��k:�U��X�K�O:��j�E*r�r�߉����eH�<6l����g�~������k'�h���X�o�Y�9����*�;j	)��H��S��1��r��1�TU*Ţ<A��.�q��@9��2vq��%b��X��G��$2�!I
��v������IU��d�����sZ���� �n�42v6�aZ����E�좮,�a���ш"����I�cN��#MȠ�H>e�W���XS�#Wj!�¬��
(HP(n�*T��
yZ�5��ĉhDs��CB�&��Vo�Z`��cl@�@����J>����):��"i�f��IT�B�f,N���z\���q����-�� �UHY9�]�ߑ���,�VYμ/�S��.�A��H��\�����1�B�*Jī5�D�k��l��HV!f�ݠ�\� ��Y������dT.�0���`DԸ,Մ�YTa��u���D�g�[WY�Y���k`b��ZNo�-I�So��v��ho׸^p��D���}+�HG�J�FW���c|��1��=�(�?i���I��%����ʰQR� �U�TjTn���iD�j�B��uv��q��3dt��#����Pa,��u}��g�`x����*8*��0Q�����;|g/<[ ��R��Sj�?&PI����D,�>����@"E&.�����54*�'=���A2���׭�H�JA�� F��Бa�#F|"[����޴�8u�3���]��Z҇4
��jDD%�);�s5z����[�	Qm/i{S��i|^�Sz�4$a� ������4IV�V�P�TDG5'7i�Lne7�	J��ŀk2���J2t��{ �MMm�����P�_Dx�$�/���̙,τ"�Yc�W�%H������x�(&3J21C����$�Q�*�!k�>�"���������?,A�(��@.���H�A�RC�x<Q%�c@d�f�	CY�7�k�Q8��\ؽ4���sG	*h�&	m�Ӎ9j,�PW� �`����Łj�E��I�#M��4�����U�J`1	Js6	��ӥb¡Ex$�-��[	#��¡+,E�0r�M��#��Et��	P��\!I�`�J `����ٜA1��xd2�˨Dq�����/�[��UJͲI��k!B��EM�(�D�cwW2
�N%$��!d���D/K��L¢͚�b�!��*Ĉ�:A��zb�B<��������ϿH�k�W��_���;���B��i�X0>�|�J�
���2c�U�|`A`�.GZ�`ǜ�����1�Eܣw�q��&d:jdԦ���j�p�-b�Y�<��Y 2)X3h&b���d�g����Fh�=8�S�>[��(ؠ �H�Sj�J��}_+�=�"��L�_��:~��*���QBP�����ԩE*��@�� �J������9�ם�R囫c�РI�2�]��]��v5G@U�	���A=b�a���Owu�ƁÌPX��A�؂\�&�k��EA!d �A������U$>��zC㋓��(ŭ`�	C��8�tn.���
J�0���	�U�qF(��k!� i1Bh��)L�b��(�s�8�f�c�ѓ8ےJR>X���Fs[�����U��u!����a0iP��b����(f�)�
���z��{�n3�%�@,&~q��7�"��@�����Wt��!�m�e]���K�@:��
����]�(��B4f7*�3n3��`�+�X`��@�5�T£�����B:9�|���P�\��Ŭ��	$E
)H$2P���JZ\5�SZ�aԍ�!J"�N�W���)hf-WHl��b��r:ʥ�W�[%���D��>��V�H(�l��"UO�_��|��vY�����{@�-�Q�0&��'2��Z��R�P�8�T���
+�у>OG��<|���뙀3�0�-ZI�ؙ�x�\�(J+6��Z
�J�q�[����J���g�FJ��&3��U@������1L�H	���{�5&�A��o[&�h��PB)"�
J��xB@X*N=��x�Y�Iʈ�t�.^�	��LbX����Qa]��1,+ $(�����H�s L�s�9�	t�ΌÚ�I2H�C���\(���� �e{���e=o�.��f#%+���ܽ4�.)���[�QuQ�w+�f����ِ�;�X��E��4�}��w��p�J���Q��"�u!�br.@ Hx�Μ�O�hU���f"��@.�����*db0@�*��l���(�A�h��ի��W��I��n7v4d|N�a
��lV��68��{���n��T	F4�W#
O��~x]�+U(��뤠�h��f5��%$^X�gƣh��H�2$$��x� �5��R���	-h�@7 KU��O.! Q$c��G0yJ\\,Q�Q׷S#�Ԡ(I:ׯ#�<�a�&<�C-���D	b" $T",H�
EQPb*0H �@"
/���gv�\�]�۹�����j"6V �nV���k8K����}(����b��2(&��6U�Mel��f�m���Mh�7��(��REC����!����LTl>�!z)r9h�R�Z���6P]ԡ���ue"��*���Q-�# >��	�.D"�hDg� �˔;��NiqdQX��>3�5\w~�S��e*� i�h �+ � ����[�m	�?����#'��!`��MTDl��F˴�1(&#�P���\����%'��z��)z` @9o��������I���Wd�imF0$H\��I�[$�f66�-�u�A0���L��i��yݎ��p0!8�X�`a�T
�f*T�ȁ5���ܧJF_�6�����?�b 1��V�hF(�H �X
���{C�tÉ�&����p\���}}�.@��8��+��Q��b��rU����^o����T�(������K^
*�P�1��K)/D�A"c��|�� �@\�0_�e�o�b�~������Z_�;�ѯ��������z�>�
"��T
��p{tO�
�� T &&�B|(��F���[��v��{ľ���KQ�p�]�&��}:X�����.�ȧ�d?3@��+����?�������q�� �pdxXug���.G�>η�˜{�W_��a��v��=ǈ����r���7������}~�Ư���L�Iv�k�����5��|�
G�v��>n��9�;��j��v��7?�v}���^���8OI��t�%�Oٙ��O����.�Z?G�x�O��v��֐>g?J,�|���Qo�~Ǽ��y�䭦���\�So��wa�����*t��}�_���?�w��{����D��9�w��?�C����\��5(f��~��K�lo�dU2!��fg<G�@���p$\��7�Gb/l�Cꡁ��P�H�]l�&��A

ZR��yQ�%��몈�C����%������Yy%wI.�NEq/hU#����'�%��v;��� ���b�&e�@�P���������_����>���������G�H��������j��� �������咷�/�Z_��/�g�<��h�p��#���?<���gf�����o�^�}m������s�[`Q)��jw��(��}S1���]Q�w�g�캌�B!��Q��>]�#V��|*\�Q��e�B�J08��f�ލ��I[,Ӭ9oF*��$!R��r��8���W5��헕�o|,z�Ou�`TO/FG��|�~�ː��w��m|_�w��϶o��y��������VqA$D^��I!�hC�v����niH�\����p�|��"|?�k=����q���?M�RK�s�ϛ�H\�!�Bx�:��GVPV5�j�,ۦ�s�Q��WwF6,Eݩ+��bQ5�;��0:�'p�!����l�S�\��*(֋b�-�,�ՌF���	�D�hKD�YZ����=������#�"�z�9��,LΖ��iI^Y��a(8��L���L�d�/����>'l�RV����$s&Fd�@�2ϗ�?"0�a:ˀVm���C�@0�	aR5 Uq���e>Y�"�aI"Hn |Y
cd��2y��I�)Er�,�;�� ������k�+{�W�͊E �ޛ�wD�.�&\utRe�u�Bbƻ�˻��խk6ש�BJ�@� &$UņEp��#���WLI$�s�r�Gu�նֲ��'��M݂����ww#%Ӗ�:sUK��9�ܔ�9\��ۥ�����SZHg9\���\��E����&"0�1�b)#���#���B`�f 9�h G}:ͩ��`bć��Ő@%O�����ٺ� ���-��B��ȶ��*�cX±����`���4)��*Ѱ�n�Ƹʰ� a����b��*Km�~K`�i ���hu7&��f�Y�g�"������5j�k�_%��(��Q��J��Q""�,E $V(� �e�� ���*��"����8n�:\���c a$\DʕU2��?>��E%�g�pYGՉih��)�i��j�2�>��TX�k7��<�4�`v�̖������=v��wu7v��5�y$��WL�Tn�2�!�f�C6̖h��H�0@��,ۑ����Q�ݬ��?4F�5KE�lJ�J�PO�nhK�l
��T
�Wa�&:-��]lp��:o���\�y(�! Q�/"	*����z"� 	+��B	�LGB�!s.�Ql�W�U��\tR��&Hc«�V&�� 
�2$�<�^y ���3w)s�G.c��� ����|�>�:yv �@��!)����p��b�a�\ M03$0�@�! T����	�M�>6g�)��u��z=��-/Ȍ�#&����dWId$ N䈴b�%��j(�B!%�<[dr�, I�S2��3l�IT]T���� ǝ�2�V���W5�Z6�k{��"T�ET$��(@&� �dAs�ـȒ$�D�*�³"�q���H_�A#���S%L�qN<��׌uс��c�>_U�>�b� �>y�j��
ǘk7��WϹO�xCdv(f���`H�|B;Y�i��E�'5���7���h�y�Ph����]6Phj�Rmg�|��������M��K��Yݻ;�(1��Y��Q01$�3i�4���Y6	�U$�\	�S)&�4ɦI4�i� D�8�fRN$�Rn���ԋQ�5
�Qd�,�4�4h �fd�ߧ~��X��ɮ}Ld�A*�2X�be�]7�i&���W:���` ե(	��4,
�\4�J���#O�/�ծ|4�y�V� @�-�(� ��0jL*��P�uóG]"ݾj���F�I��Z5��V�ZѵV�XڱUj�����X�m��hō��r-�W(�A�ޙ���~���}��%$�{����Lj+�;���d(�F߫~s���ҬljCh����k���Ȣ5$j *��F(
0@�BFE_�l�AC9�Q'������.�q�d�>y^�G65ZƷ5��7-����2*�7�wg�� `����"n_oh�D�llIQ6����_�a~���� ��w,�xt���e@BA$D$����( ���^�Y.H�~j��@�0��g��6�ǌh.���P����f�(�����$!$����>�������8ZNUWy�x�~�<|G��?��� d"v��}	<O���[���K������i퀰�@�oz:���1�|��ip*c��m�]uWp����<q�-�%b�}���X�P�^.�Hc�2�-tJ���V^,	�F!2�jJ����6�<IĞO�L�������
�����A#�|m��jw�DɊ�b%a�� �_ ��@6F��*�j����	�Q�HW�|�3�Ǻ��f &8>h���p��"GV��J�'�Ao����E����F�N��n�\Nߧ�Ob;.�(�s�5�SW�T;4@4����F՘!��6aq�x�����m������I�<(r�V nX��`}n��A/�>W�~b��∇!�"��/��=�C137��Pz����Ĺr~��3?�zFp��z��{}���=�ӀՇ���쿺p��9�U5T�?��2�a D�Uh)��{Α�{@����vR )tQ�a��%��~��-�啚�U�^�lv��D���lyB��C��69���Y6&�P� x��
5��oh�eΧ��ow����hp��m�1�I!yćpq�c"�S�Ѻ���:������\���v��"��	�N9�=�Q�b�A$DI��=���T@�A��@N��2��2��<*��"�+�(��;��	�K�t�t`>wg��P7o�1b}W�~иz�yH!�D��H����8���)���f��w^{�/j������y��:i1�^	S�	J�� ��ᔺ#���,`4t6��(/_o�-�<yJv�"W���#�7�"��"%D�$b*,[R�SH�&�$�SH@F @�$k_Wol�_��G�H ��z�=:fwr�WHy�RW@��� ����+.���bҡL��EM@٠�=��@�*	r�j���	fL�U@����ޕhhF���P2� �x%/�s!��5	!"b%���5{�ֽ(�\�@ DK@`��V�0P�`b,�X$�q���>�������7��Y4��l��J��|K<w4��{�Kv�b���B���R�E���@9@����S@�F�(D��h�n,�"�@w ��gyHH�� �Ы�/\Cl�d���Ev����}���ߧ}��A0E�I���`Ŷ�0�3 �-������]���V*9"*��t�j�������\H��dى�28(��A��
��� bS-wS:�2���lAD��g���@�FA�C�D��6o�J������}|
#TX
��Q� 5��yp���@�2 ��7mJm�Z���������~���j$���I4$���wLIM"%�M@Ыj�wWl�	#%nɪ��(�`�L�ӈD�^0���r� ���3�x�>P��W83s����b*P���T�Dȹ�d}P@�Di���!H��
.�P.YǇ�XE- �P�V� ��2��/��Dtˈ��q�BHFe!�"���ōLS��q��m�JI(j4��2�@�K\�~ρK�TQmT�%TQ@�� ���%�W��2ňj��;�� ��UP7�u���&�e.� <pȁ�W���/�dd
�b�7��J{�C(TPg����3f��a2��GI!	P�I!�� ���K��+�AsU ���fFA���4�DuQU0A��.�f*`�!��1��GP�������������H�-��j��H5�&�G�����d��,MU���_����� ��ǹ�D�(ݡV�B�@�)�Zׇ�(MJDC0"��0)q"�\�zO��'R�jg��[�lT ����`�ˤĐ�ᱍKJ�!$�h�Z!j��m���[�F� �Jc��P�wX�6s�&]����7)wS�q�b���p�4Ta6���+����-F)���!$!!@��x�bZբ�u�a,e���r���Qj"cע�];����;�n�"@��H��1$5�A5��Ԕ�2�nA� h5w
���5��cZ*<�T�,<�f-�Q�Sr�g!xC�!.Db�PǑ=*��������?G�M���u��U�.u��t�!ׅ���?v�"$��� v�5ae��;����\dA<gH�E/�b$Ѱ`�@��	p*q~r�����!�T�^$��9��|2�P�L�@ģ�*��.��h4 %cB�(M�N�0AĬ����2O��@��x�y�Cf�uۀӅg GD(s�n�Է��F��A�c��_�>�&��BI�?y�) "#	iV�/��"e# ���� ^\"�T0/�F��O����#T,� �	�DlX����^���)�10D,HX�	`t���aE���* ^A"�
<:�� ���J�~�Q���������4tگ��#��k��NgLj���RDC�b�7cn�jpa�� ;�8ts�^.�"j9,�x;��Px��b�}�i�C���<�u��N"���]P���k��q��3M� �m���������4jY��ơl���#R�l��Qne\L@o(n�	�z7I:��P�B���˝'���xr2c4^���$F�'TBM��B�YI`�N�@G���pA��L��P*�TQ@Ә�B��Ɔ�DL nP��Q,"�r�Ү�*:�U)P��i�H^���9K�گ�q���.�sF�܅	�hĮp �@�D �  *�D
Ԛ`MN�(��(E0�3��F�T��/�,I|UJ"e�t(0X�e���������F��ۥ�iFԶ CT�i�����kZBZ�rg���f��j�2YM�|ұ�Qj�z��  P�(�`�&�!�&耙,��ż����b�� i��p9�~h=�1��r�(�DAc\���PB��<��r!�iǹ3�HNP0�^$GNf�
\&!6�	��.� q#Y�"�I�Eհ4P���$�����:G���9���P�i�Vx;؂j���*&�72D�z &+Ɨ"�~��|�Ed@�~�e
��n�$�6-@�>;fK�PCDH~LJ�~�z^~1,'
�4@�:�t�0x����� �"	"
����qv�H����M�I��
���m�TW�=�;z ^k���k_�1(+���X���r5!��y��=X��$<�'f�!!&L���=:pjR�B@;�q�I }��$���PE�,	P����hZ���y�;@h�!̩_8�H�/ido��w�,)�7���t����A *���%�d����K��X�޼�@o��'���) �3S�n7ER��j,��~Cf�X ���RX��&��X}LP����x^��PK����}&����|�\���q�_�����ɟ�v��{.�v��K~�^���X�݊����vO����v"��FEEg�=�e[ q��'^VV�|����8�Y��y칟c}�a�ω��Ǐ��frv���*[+��o��_�k�,���¿r�&�G�m�������4���o����ﾏ|L���>�$r����C�Xf�$_8ؘ@rNPh~�W�L'��,���Z�����u�<[=5�Y���"�&�1z���~������W��o���7�_��i�;�?�������x�#~�W��ݏ�������y.�z���{>�������w���g����#��������oa'����Ȯ�2�o�yG�l\�kC�h>Qi�.d�ԂIo�?���<K��s�O�J�{}��q���,qJ���~���nz���z�o�<�E�~���ʫ>P�G��Οc	���H�����h_��}����؟7��}���?������/�O�{����c������T1u��|K������g�m���Y��o�H��Q�w�����c�t�t����!=�Ú�*�/��?�?_�+���y/�߰+�{�+�׋�i�;}��	�
�=��|��a#$O��/��m�1�VH[����ӧ��K�I�Oa��M�u�^[i�����p�O/�t]G)�z[������p^���߇缷aq�O���feFn��(�у��㢻J��9�M���v�f�adr�ٱ3'�����?��Г�k|�J��bD�}���2m�t>g������w�?��.�o���^��{ӟ����:���6���Tt�_��w����5i�y�_V��?U��!V��?����_t���~�ɩ7��>-�a�����o���o�=�|�����/��:/����}�?����}���0�~��gg�Z��P�������v"p�i�������t��:V?�O�!�//���%�c/3���x.!إ8Q�mWo�6wNZV�!��u��T����F��R}^��I���^��}�I����?���~����`x@$d\���ޥ��!�F!�7_c�\z�� @!��5��.��v�6���ja1�h�7Sk�֟�s����?�ԅ�g�k�_bY �(�������=�]��D9�s3U��7���ܼ�1�>7���t9��j}6K��#���<T޹O��o����I��a���z���?��_=�=O��Fܳ��������&���_A��7����7wE����{O�_��+������8{����?��H�^x^^_�{����_��Wm�}�ݿ+�j�?q�y��{���}U��w���g���~go��y]���]���.c���XF~g��/�[������?O����s�~Z2|e��-�C�����?��!���k=D%��+�?'���z��E?7����j�������sM���W����;����L>����Yz9��p��?��s����_��hN7�/�~Ӫ_���������'�W��.f~�8y��O���_��I'���a�[�����.����#������!�O���[�=�O�����H����#�S�*��������s�?��������{��n���?��8|}���þ����n��+�#�˾�����J��|�W�;��~�j����}����{ϓ���o�������_НET����o����_q ����� �,���Q�~o��+��'��<�S��K���W��Y�=/��#��>�H����o<�r������T�o����s?�Oڷ��������}�xQ�y�����Wꭄ.{��S�|��?��3�����_����;���>b#��ǳe_��'x�ހ���C�5�������N�W��E�&����7��v�g��o�m��9�3�p^�����d����G���۫���}u�7��)f1l��;���F�7Җ��.����ߒ��n9���7t�-�=#���qf{���7���x]�������������\��?�i,A@��i4�'a����������� �
*�@C��=l�x����Hj��,��)"v��[ZR�!za�B�Jk��c�Td2�4VUB*��Rc���YM���R�|/���r�8�+, �r���r���мB�DW�7E��|�B��Dm���U��t����)|C�$^ �(Qt�L�t�^c���$E/�}��oM�~��e�o[��u�������=@�r;��#�q��/o����E2r;/!�%�`��w�}L(KN�P~6�P��$��K�Đ�C�(S�P��?2����n��R{�=����T	6�N��}�c�)�y�)$d���iOĐ���)hDR������/�|�ݒH��.>�A�I�(!�� �)i��'i���i@w�aqU�
����'�oh��0-�%����\.8|��q�{4�~�t��ԡ8U�G�`�����y�=O(Ui����:�/>���?�r<�$?�w���q�=�̝>��\��q��B�,}��93�.8�"��'�"s�>P|D���B��yP).:�������!�y��ϯ	�\��z ��K�L1O����н�,*�q^X ��{õ��\�$)9����.=A9���^>���^��}��B�Q$uGfI$��I���
�% 3ȕG��"$�@(""��E $V1T��"��� ����V]r|��!p�"� �X�@" "@"�T����e.@A@ ~��!KaVE$D ���?l��oE	��'����qz�B��VUJ��m�mJ�ڊ�B"E�W������ +h����2�B�(����\
2*� �ه��B�.A�0V5�jj�R�-Ml��TD�1ǫ��2�DF@�؝�� H�
� #�/�G$]�\�N4r�Q�J�!��f��D�E�1;ʱ��U a��K�ݳ{_s�:�i;��l�|�G�=����4��޽�,ג��:{snν��o��6���rFN�ɀ� 	�MkZZs�N�&����f�^Mt� C�'nW4w���\��ۑ�59S�P���.&��U��L���qz��]�{�v,�؎�۸��2a�%��,�&U����y3P9b
^�J�ԭ5Sm-��U�l��f�ڦ��J��kKHP���p~��M��m	��˜t��V�����?�ڈ�G���ݚ?�1J*�_���,q�V��]
Y�\^����**�iV
�a�e*���%e��
�F,L1j��.��V���0��Ԍ����x���ޮt�]����U��)N��Y4D��ڱ�!Y����NTr�+������0C��E@ �8�c��˳-��,َϜ�r\�V`v���Ѝ-������D6�'&cGl��&�mZ?9Ҹ\F�e�v�/GH�Kl⸜6��q�R&a��+;�G���B��bp}ﵱ5�Y�6�m������u�O��3��Y�n��4ys��K?W1��]oH�魭��՞E���.���ի���+i*.�$�_M"��������J�F�sN&�''E��-���!5����i��W�x��8f݊���N�|q��I7��t��D"� k�={����{N��W�����w���Е|?̭���R3�>z�N�2�'��YCm��a
����zc��/�9�(�?E�aU5�F�lNz�yj��[q�h4�F�Zs�j'>��)J���:�;b\�A6t,�qX-wU|sq=��#7q�)I𱽷|�-V��2������U��.�G���.��k������D^҆��S7�k�H��q���ه5~�Ƽ⳴7�8���������:88ә��<ar�SK�eMy���*�h�G����ۤ�{�!��E�F�W��ӧ�?�� ��PbAE�� !����m������]�q��n��O�/w�a��a��ee���*5�^�^H�כ��cn��a�^`�_Md�bzZ�aM7Y�{�m[>9�Y����?Pc�9~+��=��Ƃ�q����T��rW1���ezmH@BWb��w�oZ�.jm�u��t�|v�]��S�nݫ�騆e[�3�ߦ7�+�՜�\_~��Aߛ�G�$׃��Ӹu6��b�u����#߭\;5c\t�k�y}!~uټ.�#��z]�I��x����Ӯ���pc�kN�R��[�s�=7�\��H_�y��~ԥy=1Jw�e掓b]��/��\�|u�v�^�ӊ��������}<j�x3:ej����NM1�X�����~B\�
`��<��k-�%�����E�%�b�@�"�H Ab,"�H� `�@u����l<��Ec׿��? ���������Uo-i�Wߏ�ph !�zڱ�O�}������G��>4����!E��zyvk�f��������]zz��TX��jwc���s�a��^k�:���6gB�9��������������\zO�^:Y�����kq���^��am�)��]�F=#o1�1�k׫�{_�]o�/�yw����U��i�������@j���m`mӨ��{�]��璘~ԻO�z���o�N�m�3On�5�z=��i�=WNk�V{��>=׌֒��>6��;�����s�ݽw�i��k������펜�1�g������j���q�.ݷ�5�u�{�כ�˯_'�)���0����=� ��'Q�g�_Ou�m�m�=�*�;�֜׾�i�ׯ�Շ����nޏ�|���}�y������S[k����4��t9߫�� ������ �
" � �Mm�lu�z{z�3��Wc�:��"IE�6'I��W�bBcň��lҋXi
�wpUU;_S�[�O����==,���^Xu�:P���/���1�i�����&H�(*�0���Ӣ8L�*���g�Oe��}a9�4�IC�L!eƏ��9�D"�0х&�&YL��w���;�s��K����l��Y�h��a�'�m��c�&��6҅��K@Ƥ�K��'��ȃ��2�h�8��,s�}7���_.���|��Y{|.}�> ��v����{�~�	�JL��
�ێ�(�&�i��U�.lB�����=��w���*�juvt�h�{��k�{��F����;������6��tھ���ۧ��Q���i��߼)�W|p����0#K*��
��8�n8j���e��� U�c2th�$��J�<�a��Pn2d.����Ɩ��4���8����I�M<�����}�N�q����M��S�w�v_j>���wϹ�I�a��{q���w��vV8�_dO�h����_��0� D ����  ��O���IRɮ�h�Ů�Z��ud�%�L��2X(��DO�5�k=�G&�yaB*w�'�(�;(�H�&��@�4�Ө0X�M�n�턐0A��u�J'���\��/U�����{W��]�u�]��릚����~{�>���o7���H򺮰��TJ�����s����x$s�<ͣ�ΐH&���lK�\P# �&K���7��IW$�m��r
�cC��٫NY��5ǂ��	\�ɳ8LC:�1�<�0���1�,,j�������HOTԁ	"@����,봳��4�O��<aJ�3/��A���������]ea����2Ǆȝnh�l�S8�
H����3���$;�)"�������a�0d��F�� H��j��2����>;����JO���=���}i��ǟ��5�צԧ����!O���1}�>����~���_���u𴮛|6�{���%�3�y�~-��H����>�O�4e����|���V�z��|��H��Z�O�.^���m҂q�ڕ�k��Q�o^�R�Y�K,�K�ɍL3 8� �F�pi� �B1��B��Ԭ��Ӽ������ã���M������+��$I$�O��7T7���$�! *�7t���a�kw}�����l�@�@�#_焋
�H�%�
�I�] �\���
��� �,�����͎��W"v5y�����)b��Ė�ޤ@�vzZ�����@�b�Y��-障i 	ȩ��-TȔx�}��7�r9߅���TVf5TQ���P�r����<��{r@(��<�T�A<�b�\�1�HXN�-;0�sR҆� h �x�T��
BgLeׅxk���(sOh��t"�#D��4sN��BB!H��#Z�&@r
b�l�F1U�Bn���,����K`��U��R��Ϡ�Ȝ�UL���2D��~��	XՈ5�2`@�4قr�8�?-fN9G�wT
A��Dbu���z]~!U�96_9�f �X�@����d��~g����X��.󯱦��H�Ϯ�0U�{�{�~l7^T��aU��u������z��h���0
��+\@`@Y��QD�Tf����5�N��V R�q�J*FR��a��$�D��rxb��Ve!p�b ��	:�IO;~���cbEp��)B���q��r�����<�2���JOlȓY%�8��)�������H�y�%4��*2�����1j�~~L�ݛS�?`���� �@ ,kf�ږ�TՖ����$E�V(DX#"1V" <���.��*���]���R�{�&�F&�N̯ �;	e.���\��~��%X��k�^�
�6A���l(��$cB�P�6�_5����N��8�h@��h�&`L�	�g&��
�:dڦ+u/=�T�\��	+pӅD���ǅ8d��㒒��\��'2�	!z#��Z�H��s;��oq��h���� 8�EN\b�9Kgą�/QD��)�v!��X� �P
�����-C��SV�����Q.�㸶�A��it�$p&R�Zry#��C8*�YKE#ν�d����[�=.�:/+HjBۤ�h�Ȍ�423�Ϣ�-:��MjC6��� xgz�I�����ݘfH�AY�d��%����
#�tMJ�)[.-x�0PKFZ������ME�PL��z�!�׋0D�F�,�LQ�zL�	��B��޺q�0�8�g�Q�@���{��I�8
VF]4jHKp� 8J��4Y��i��P�* �$0�D3�rzfI��(�
���Kt���jS���YWF�D����}�Qz�Zh�.I:&x�˞�����%E�a�X�$c&BL�4$آo
�qz�&\��E��G�fH�1���n:j�-B�)b���ZV X���#�`�0JFذKd:�Xs�P`+1����] �3cZ1�3������t+�89�-<[���|��F��P""� �2(#x�n�ޫa��w>�i�����n5�{�����K[�[_��<�/��L�j-)��i�]�53��x�,���,�F!���f�WF���!�Q��������+"RVN#������02d4!:[fv0�d�Y�0#R��1Uڵ�l�|Є!Rr�^�ybF@�ϱ�y+#�f��_
j�DoMT��L(X�\+�����pVd�AJԌ��P���j &s)�\B0��*1"�"�K�Pe��rY$�J���b�b�E 켋���Cw��Դ� �Sl8BID
I�3�"b& 6"K	 �m�S
D��+��K5;�����dD�66X�@$�)U��ۥN*iZ놕�>$�fT2p�`!��\�fDT�q�V�%$����
4v**A�r�rs�-�H�����`�OA��o�=ᜐ=����O$U;@�崚I��܂J$^�1�	=����:�p�㯀��,��|7���Z����&�1AS�T���n���}�G":ƈ��Ș�3�X�ߊvUVN.#^bJ$VG$ %ٝ��!�K�Ȕ�:\���O��L�'�\���S,q ��H���2>r�c�ԨW�	��Z��]m<�O����bB�Y�L�.�FQ&��E�U��a� 0$�e��V`�䞷���&]Z�"
MZ@��:��:I" �6 �"�pȐ,7<���5�\��J����Ē���nx��`N�H$�};�&�7sC2���8vޖ���k*7��!�����]�)2�@g+�)�e�Bjp�G~ӫ���Ķ�m%E�?�y�`��� �@�� 'e������5�C@G �8R�<�D?J�8C8���-6�R�?*/�D5�N)���&$�^�T	Y0�Q6�\B�8-�p�bx�ޗ�,�$�Sޢ���F`����ϩ"	C�=�ͥJ%��%����7(eߑ�P��^T0b��mAm7x�2�.�x<�`�7�RB��RDF�� D���?x
�v���!����$�j�`�4�� g�E�()���K �8�`u]YSO�`'�c`<X�,�nm�U�<C0+�c�ζ��x-�[����茈j��z�v�&.YUW���8�T�յ��V5A[��7
�b�@mwa���ִG�;dFԓ�h�.�G�1��RXD%`h�-x�R�D�?0==J���\�W��e���"j�zSHq�mM7�����'����]�ύ���z������F��N"�e�x��U�L�:] f�%�R�p��]F�@�a�d'_	;��x"X�m��ؕRі<��W��%�Yy`����6�$�Kk顅0�@uf����"����p*�Q���N���&��P=Ӝ�a٣�a�eQ�l �#��;D��:Xr�*�dr��l�����\`�AuG�{�d��#�`��X��(�I| %���Cfo�%31����%	�%k�N��:!����͸�xΕ���D��� �83!�Ә���ԣl��f�qg�K|�Ĭ����"�,R�3�+��:ã�]�l8�D�95�QV���X%ԁ�7��aj�l��)^p�\�̵/TV�7�U��L���T�/�p�V��w���v~�n۶��-moڝ���~���h}>R����d�x������BA��P��Fߗ%����bd��[�[X��mmZ6��6�ۼ�⻵���B���ì�nUw]�t�Uun&�:�%��M��j�[�kl`�U b���Z�V�6���fD�&@�)%$��j�(���)hā��F4l��+(زĲ�kB1���[k�y��2ܱj�b4`�`5lZ�����D[��j�E�+��j+��\��TZ�˻mD1���mTmFѴTo��չh��ʍ��r�r��Q�Z�W+�r�� T%I�ȡ�9�}�>7���7��~�����>O�����߽��\������C�������_a�?������������������y���������?��?�s=�v������:*A�dR���"�h�LD����F�5X��%l��[Zɴh�b�5��Qmhډ6�(�ʵ��j���VA6�k�Dmh�6�VA�f���D�ʂ(J�V�-V�V6�m��mh�@�[b֤aP)��P؍6�Z*ѣR[lm�[cj�kZ�F����Uk��kV5m��j+cZ������QU�-Q�����Ũ�ѭ��ѵm�Qmj�Q�[��j��F�b�صcUcmb���Q�Q�5cZ��F�ѭ��klZ֍�F����"B��A���P* !IX(Z� Y�縏�{������7)�����N��1�����?������ˮ���k��7��o/����o�z~���G���<_�k}�a��{�[��]�o�o�{oe���?���w~�O��)�;��5[��,Z-Le��$dYL��" H�2AF0��1�`1�(BL�ifa`�	"b2	��ً�b� �E��3$�21��LI�&b�Qc$R&%L�$,�`%30���̒�H�AK2�R�L#")Bf�L��B,$�L"1#2b�ĔBDBRH%�H�HI2@�$�I1�(�%e&� ����2D҈"��J%6$�!��4�1RP�)���JBZP�E%�I �,,J�&�$&�i�3�"�hdd���SH�1�dē4d̦ɓ"�"@�4kLi(� $H Đ�i3I�3���Id����$�S1��dH#4҄B2@ �0(���$��ģM��531��cd��4�@ j��#���g��?ץ�;�������Q�j�o��<���?o��>�t��W��_7�~���㻿C� P�+p����Wk����ۼ����^Ǹ���ߏ���3~���~Ϝ�_O��m��}.۶=Q����w��?��u�}U��?�v^����;k�'��m��;�v���ޣi��ߊ�;�v^~?[��߽��<��"�)_�*?�(4�] �l�@��]��=����DQe��4���1^��:��O�~C���L1�B�K�?����ACrNfMw���	����|���l�F�&#���2��%��C���K����;���4���¯�+W�8C8�������I�)�L�<
uJ[$g�����H.��L��`�r��&�)�1+sVW,��`$Ջ�/4B�:im�*�E�T���WL�I�H��N�����j�����vN��怜�v�Q��}���\���Ab��U��4��H��K�C���(�dB�9�n����cNmUZṇURQ�T�KU�c��%8;�:�%�F�g����>5�;-���b�$����4kS<e�f%ʶh�ED�^<v���`Ge*ӆx���'���A��֡(�a>Vr���I���9Nз�_2I�T���������aA$i,�-��tw�9�m�>-[X<.���\� k8���D�K~�"JbMM0>H�s�5&�|8�z(� @f����kH̺"�d�CEU���o�ܓ�B4g#�#*&5CVM6�)��p#`���u�q���9�-���i�E�\���x^W]�HwCR�3�� #(UΪ�e��e�e�a�	�ZD�f��������;���<����1���/̸oι��ͤ�ċQ��8�9a��X��(c��JCDS�%�
BA�"�;�P��%�"�X�5�kXy�$��u���P+���1�GV�PN@�J|"G4y?�B� ��朡��̈�Fj.�w��s���|�j?n�w�V���%��m%���@�L���cR���1���y y yr��;���� ��C�A_��O�i��=��#R��@au��"�,T27��10���0���F�'���}Z��'���8�ń��R�Rd�h��Q�n����SSʉ|�.j*����K��;�-B�@�\!�.�(d�U��c�$��Ҥ�������r5��Z���m�m�66����^�דڭ�i�x���FV0n�
���� ����/UU���*�T EZ�����`(��(��A�- UB������� �T�&lP�-2ZP��mI ��-A��\�TKE3*�1�*�\V��_E��p���A�B�KE�q��R�|Sn��j���\1�$�� +PH�)PD$D�@�(��Bd�b 7E$A<1T7o�y�:��A�2��V��V��&#���e5��_��?�_������������������������������������B��a�@�(v�    �Z�W�A:�        �             �             �   7w�@ I��@6ƀ2R(�P���          �(�.
(�ܹ�tn   w |p����   }�sI����(R�	� ����   �[� D�zM�,`<   �4�rNP  �h�   p 8� �   ���  ^    ��޽    O�                                   ��H  ;�   ��9�  w���g�>�KF�   �()Q��Q%!*$��e*H�M�   :R�BQ@H�P� 
�E;���j�@
 � ��70   :��am��8�A���	�)��͆�m(ш�f�m�II����a�Q(`J����v�ܸϖp�v^� ���q�xy�  t ��*�` ` �!QB�s� Ѹ@    ����
��     � �@��4��F4f��&��	�15�2=	�j{Q������=MS�OE=�~��SFM�?�H�Ğ�J4 d  L�	��m5M��~����Ci<���x��M�O4)�1��̧���'�Q��ȧ�&�z@ SCM ڍ�A� &�d�CAR�R�&ѡSC@d���M �&�4  ��h �     �       	4��DI�&4�z�?S#@#5�L�F�P��&F4i����di�4ɣ hhɠa4� �h� ���@@�bd���ɢ��e<��OSOQ�='��@�@�4������mF�6PPd�4d��hzj�� F����������	�	�3ɦMA�����	�	�`i�ɑ��i�hɦS?M40FL�2�i�2dMS��P�E��%م/IS0�_����m77.5�Msi�hɮm5K�8t�q}���`���3.��Oڟz���]w�5�m~=�s"s.!���ЊsR�q��>V�IK�DD�	����ٯ9'�q�E��9vT�LɘW=�u�<ϝ�v�����҂	����UJ�S7�0J�v�f�+�|��g�~{�k���jL(��%yL�z�fUK�G�jAN��~��/������"V��O���`[������Ϊl0d
Ԧ�"@"*�_�f�I�AEO�YC��PDX�f�G����U���\�m�ٚF2,��~��d�R[`$�H���~�3AARҫ�KEV8�SB�1DDk*�ʌݵ�UP6���(����s]LER�'��c��2���6�Ժ�DQg7(�EH��ē�h�����Д|��|�W`��t�UK�*�t@Ǣ��Ԇݐ1߽����2�H�?���6����m����띡�1Ke���0��_Sz�Ҳ�QE]��eˏ�ڦR�Z:�m;
�R�� �m
�L;U'˫JrJեB5)^����I��T�O����O�����G���.&��/����*��������w*���1TjҴm�S2@�$�lаU2^�ZU�\���g:{ٟx&& `��� ��	!��$�^'��)mjٴ�ʖ�~8g�$�>F �>��܆�,]O�ɰ�$������4�����/;�!�M��� @؀�@�O���׿Iߋ1��@fڌ�;��g�W����B>�-k8v{��N3���ٹ��j�<��k!Q�����W5�i;Ύ�`g��J�!�����@�B��+Mj���"Ȓ4�z�o��?A�+�k����lUx�	�3��P
oΛުdTs,��Ҫ����5�-Q��ˇ�z~3�����z���)U.�����]��V�TP�ֲ�!ȥ�m��V�f�-2�-�3�R���;�*�R�*(��SQiYǘ%�DD��m��1>��b��a�,�um��mSYq�&0�h�/�s����"[�]���:�+�c{ώ&2�S��L�Uc�G�ܾ�W�.%*�fcY�N�͖�h�"V���߮�X��^�1֣��|nncW3l]i�]g��;�R\�����n�[[w%T˻���H_��,��(�*�ޭ�۴��0��
�(�J�JRUj +��~�"�X��r1B�/��0=�4r���\pX[��0c11j8�3.���I�i��	����[d��U�D �s�f����t����}�O��?�e�}�oO��6�K"�k�� �f���?����:m���z��ʠ*��S�{�N$�qE�T��TRPo%�1�36���E���f&�w���츩����R�#Z�B�K�1V�Ma�2��Q�"���fPJ�[����nmL���55�a���6ܯ�(�
l���Z&��2�Q���ؖ���.�{3%W����)�fR�+i]�e�6ˍ�VԢ��EUa%�hl��.ڊ�%TX���"�eE�*�$Lj
1��c7`T\�čܗ3kd�4�Rݭ�T]u57r�i�Eo��� Qbȉ|���ۋ���ʕ1���2+���f���C'��5���sΧ��]�nfQˍ�ˎu��TF�5��/m�̓-�ۘ�b�Q�1ͣ��.�HHC�rw*�2���W]A��(�!�d�땦5���wn��6�b[s�ݳ1�(c�*����j�Rҡe��n&ikr�q�T�7sjk�ڶaEwAO�]��2��ۆ����us�s�U���]w=�g�U5�o_>��km18����`ݦ9U]W��=���˙��m��a]��.��s�&�dw���Q����Ki�=�h89��jV��3(����\��TnaF]ʹ�%8V�ݦ737&\ǫ�;3�����nU˻(��(�Y��m˙�9|��|����GOn���+�=��m�Om]�V黨�R�+�Gr�u+���n8R٢�#��:���҃�2�]�0҉��qLLN��/J������543z��^���m�k�p�z�ʥ�F�&e��)�V\�aJ�o���9�"��]z�f��7J[v�yͶ�ۙٷk+�vB�[�s3�!	$��۽��v�Hڊ�Vh�mM��r����b��S�b�QF��m[[Y�m���dmV͓͌e�b��6����l_?�fj̶m�#"M����Y�Rؒ"��$����M���5Lɳo��౉�ZHX�#b�� ,�E�6���}���j����	����$UUm8Έ�~]E}>ɮ?�L)r���{�"�h� �h,SI�E����+@#��v��U�WewU^p+��UW%/�d0)}@*��Z�[jɯ#��J`c�]�T�Z � ��S�2,����5L���T"�1���2%ݦ� (ez,lKv�T@ Єm��i��q��z�r�|0�F'��u������_������{t��7��Yx|r�����״�?��d[�i����;�?��7�����?������Ǒ����_��o��}'�����=c鿝�s��<�λ�)��t#���?t���</ʸ��]���z�[��}�}_gf�]����{���}k�!#|_��{�o�_Y��?��96��|b�#��Ys=>w�ו̌r���2����}_�V�(6������1�7��"��>Ǖ~�����F>��+���¹y���}�"|���\�M� �u����^��k��Ϩ���}�c�~M��S�rm���;�|�f�}߭�W��s��� ��YS;��{V����}�O��M�-�澎��kwxߕ����{$|�y��lPL~|��>����E�u��9���z�W�}�_o/��?[����_rŻ��?_L���y�yx�����*����>�������ok�2��}g��^����u�\�-������ߟ�N�5�[z'd�����J>�[�<_���{���a����hI���}����tz����7�Sf��g���yt��|����7��?�}��s� >���f^,E�x�����=��n��I�$�Nz
{������Y�w�����Sq�yͯG�����g��f�Oo��e����l�ES��x9���ٳ8��-��p�v���Y�b]�CEH	�1�W�<�������? �q��8�o}����fO�j�{c�:�s�U28Y
L����{��x C�]����͹P ɫ(,l��C{�P B|�>&%�"xF�� G|>�FD!$  ���%�J�剹\�O�.�}��(R���o`p<�! ! �%?r���`pG?zP0#��><IÏ�L[�x �Ic�bB-�����N��'	O��y��-�!��4Z,���k����  v�����8�An�����\|�8R��-��R�fY{qm��  - �@� �����}I� 2�⺹�_y�Kq2)V�^���G�����]4�  ����
��kT��ú�V�9>��ݎ�gQ ! �=D��1 � z�Uo��x�x�S���9�+�\j @!�*k)�}zr����oC�	RQ�u���j�ʀ�@ �XՄ�Y������'��G�]8@꣗c�o�\��S�L;BԛX���R��@�죔���_}�;�lXO`J��O�y�!�+��g2�\� 0!B�C���	���m46�ꢞW8��ڨ��ʊ
.�AU�(�A���ez���p�؄��ԉiС����f^<RŽ�v��^�؞=���P �E�����#�����'���tA�oNA��ܸt��>L61P]<�B �-��)Z���<��꾼v ����g yt�v9�Rw�   ,p���j;(��&y��o���+�f�@ �����E�v8z����n��   �F�������-䤀�z�n�R���e�Rˎ�ی @ 1��
͗��.E�u/�3m$#cY!h�wj�]�.�>�W��� �!������-���ҷ#�Ħ��s 󍼻�hNf�BP��><�J����a� @ 	(�TKXL<<1�(�y�,| ����#;_���+�d���� ̄!Bi�5E���e�&�7��㭇���%���\֯~���B�6Fw�W3�:������;�S5��"�   XI��3:d�{f����n�De$�.IMk!a@  Z�wf=(N6�SAmK~j].��[k�+2�K�R�o��+�)�:��b�!	���2Ζ�Mt��k8nr�o��e4�Q�(@  �$�	�m�U��P{��M�:57Іm��|��G�<l���o7��  2Ǟ3v>Kƍ/��z��A.�����q��^ց @�����h��3����G ��U:��z8�{�=S���+_�`˿(	�Z<   �<g%@N(��v!]Qb��Z
��2  ��y9:����${�2�^>[b�@@�`^�n/�5�j�}P�@!1�Zה;�=U���q�{�W��L1 Bw�;Q�LFK!R����q��ͨ}��q�/� @ �ȷ6�#z���ɮ��M��LT'A�T�/n0��
���  +�[���� �B�  
@Q����;���� @��  HB��9$ �h>��'�^����Q�&�
N�4��aǯQ�c��  �9����5�:S���ヶ�  �7udm3��t�v��2�N*�}N���tO��$5�  =B�8x�ru�n����+ṯ��;� W��  �Q�yٟ.J��<��><o�]0��#��T���N� �65����	Ɏ1�;��)A~;ל��1Y�����7굩h�  E�Pn ��7�����y7�҃z�]l9L��!�  ��t4�u�6'a�e�Vnv�k��燏����H�~�9Iͻm��<
�8�6@�  kx��U��)�)�Ne���6�L@  /W�&����wa|7��#�K�J�K�W�G � � @ �/Wl�k�ґ��|xq�)aյ��s~�� �����!U��"n��� ���@�h�݋殝�JZ=��Y �d�E���ph����@!W&���C��)�hc_����������1]\B �)!,]������k��鯹��Ѐ@  b������ݸ�Z�]�A�_k+���ˀ��GS8��H=�E�Mk�J�I@��̣O�@  	�B�w��A�ݘy%t��Sg����������H��=ׯEQ������v�x�  �(on�q����^^��\�3��T� ����4��*�3��,z�%K�ם���B�t���*����B���:h�-\�����k���/��韙�  ��ֺ9̂�?|c%�|��a�S���'L_��x��� F�a�ʙ�I�!݃�n�2Jك�@!  ;���|���,`s����:��� �!BT�I���,��c����E@��[U���
��WH�)�h������8��nj�5S��f֪k�{.e�9�����mL-���1*6)h�Ԝ�ac�f�ŭ�]w*�Z�)�u�q3;ټ��Kl̵�L��iL-�R����Y�3w.���[�1�D�� 0����l�[K�Dݦx��.�{hT���9e�fz鶩)l�S��Y�U��!)���1
��rH4���P��`��5*S���[�n]ss1��0��w3����Y�6��A���wm�1���|������wS�3��DW�3;;��
&�Q*�&Ze���\놶�X+���r~�jr��J��=�p5�i�`�w*��{�7.sQu��J�:�KN}ٱ�[�15�{*l�ܕ�L���m����-����˻��6�1+�G-ML1�,AMq׭�·.v�e1���u��-�b9����qX��r���x��ܥ�b�Pݨx!�G[l���4�*�o�ιSv+�bb��3,6�Xwfm��Wv�j��r5�c)KR�f"�QU�D�k0̵��ˮjc��;��v�떨�a�����m�]������Z&��w�k�5�WKFۛh�4њm�s{Mڼ���Ab����Y��U]˓\[�aZ�W�{�v9�V�&�j[JZ�nc1�&[i�tεq�a�[r��sݹTԦ��1��*���-��w�c�嫽�����+�q���Q��:�q����0�2�ʖ�Ms�J�˾�nˌF���,�o�&ަ��U��5���K{�/S&�k9;h�Ҙ�^�71��vZ���|ܮ�m4�]+�n��/U��f	K�Zò��v��\�W�$�E1�Kje�V޺�;�S��ͭ�QV(�-��"��Qr������_'<�[Zn�t��*v����*ڪ4��;0���;(��9�m�srӻ}�0ҹ/���R����̮�NF�̷�h��tn�l�_H ����{��!��n&u��fU
�)نo\�PNBܷ�m9�sw;������,����K���j6��:��4pD�@�ј�Sψ�K�<�s��OH�ulKb^�3ٮ赕�nbTYr�v��r*6�;-ۂZ�p�LJ��+�뮮����]1\nZ�W.�.W\�z��Uy���:wU��-r�6	Zq����E�ۗ\����u51�y��8�k;1u�9���r�L3�W)U4�m�Z�%j��nZ��a��C�K�j��=��׫��=k��zB���feC�jva�nK1�	v���뭫���q͎Js�a�GfA���J�6�pjbm���w.6^̘Zr`ȣ�j,�76��S��\�y3�{Tv׹+������cbm�KJ�5�Z��n�)���k�
뙹Z�]C�v�[n�㽻�6�:�t���F\:�:�4���n��h�2���c��r¤�6�f��5KL��SiÂ]�h�cU����휕�	���m�(��O'a�$�|_8'2� �{2��Bd�]�s�^	�g��������z��@{kw��E/�	!����q��������[L=�]��6�0�l�ܩL�Q��Q�u��֢.Ӻ��캃��ۍ(�nXm��ٻ���{�z���C�D�w3+��+5�Z�j��G�9f�E[��}�	��z�fk�<�ӷ�Q��˅��wf;Cm7[�kWɘ����J����.�_Xrc9�ögV�u:qUK醼�.睦���M�^��f;����ǚ�9�a�̢3-�*ڥ�܆\�llS\C)E9ܵ׭-���KS��]-;;5*;pņfy�]��m����eB�K�ni����ȮQcTˇZ_N7T�j�OS=�Ħ%�0S8>�Ǉ������:�g5D1(%FҴ��+��enXn]�\S�9�e�v��-�\99\Ԧer���={/&w�r=m)mX��*��:j�b�m=��N�R��c�ޯSS�v�n�NpT9+*9����7(�KZ����TԺ�Z�R����b���On*[e-˘gnw���q�����+y
���֬�}��c-�DmQE��3s#��e�S^��v]�\�Ɨnb�[c}��=%��;ۺ[U����Q��F�r���=2Sm����,�U�\��h�존��fnڝ�ɧR�l"��U-R�S�as�;ng9F��|ۏ̢=i+.�r���gf`�f>��{�Ond��]vV�K�33�rnU$�f&)��q�ĥ)K^��q�,�����&u/v�׌��ىG-�7)\��[fT�[+�w)��fS��SKf�����ݻ����������ڏ�w�.�yr�w�k�)+�y��s�M��wi�:�KU�Tf1�U��UƯ�ջ�V�G���[]����v�7�B��71U_5�V��c�쩖�+��J�s+���2��s;8�x5.S�rk�3�Qwf#��1��|�q��wwfy�w��K{�ŵ{)l�ku�jvC7
��z�2�ĵ)]��
����L��Lf-��`��{rw\��k�X�{���*o��m,�s�o���]w0}�+�T�+\)��irʍV��3DFe�]b�Je-a]��4q��[mwn�]�7�n����³v���{/!v�8"�T��3�K�h��fЮ:�:Yv���ܳ5+��)�-E2�q�`33v��wv��b9�U9�t�Ƨ�Kj�k�u1�|��\DIK�˶����Pz�(�\US^ww3�f��*�
b�n�S�]Q����{*b�)w&mV[W�W}a����T��Yaqi��־LN������'Z�Y�J��qLj��}v��=��\rұ�q�܋��9�n^w
�����8�/�*�0��y�r�rUq��D�̬r�=�᪜�..va��kY��1Xi���g[�L�qZ(��.�Ki���Z�M���f������.�r�4b'u{p���5c\LC-��4����;���q����X[k.��v�\�Xu9�˻X��q��v����mb���e�LJ��2�,P�T��K�V�1\p�fg�f྇�����֕ln[׻z�uκ�Z�z�1M��a\�Q�7w�G�b��nn�z�b�K�s.732�R�m��f:�n���7p�R�iA�k.Y�Ev�+m��3z�|{p�e�.]��Y^��KiDV������fӚ�R̯i���N�\�r��K�Du��F�`�*dys��3C��jWR�a�+Z(����mθ��2�����y=n6�;��l0QL�F��L\]�ܸĭ1m�k)^����s
�JQ�KV޵�h��Q=nJ-��-q닙�w6�}��w�4�ۑi�p�rX��˖�����E[sj��ج�\k1�˗-�ܧev���'7k���s.��FT6��+EQˆ-UY[-�B�S����:7n[3c�JT�W��v�lb��\���&c+�r���
�:YmYh�"���n�<�6d�j�]�6aG(u��w�1��]W\jm�0�I�jM�Ħ��u3����0���mǌ͢U��h�&�n�L�ͷh��c����u̹�e*��[P�XW6�nY��-��:�o���u��Jfd�)J�cM��ڈ^��^���-�*��n�ULqDťq�ˉ�ۘ��n�v��e˅�2�-^pTD��nu��9����jV�o[��Y�Z�/����_6aiF�(���1�ے�h�2�ULێ�ak�e^N�im;sU4�����陘�VշneRUJޡXm,5mX�R[LLUy��Vw���P���[o�7nvY�y�Nh�m�f�AZQ�[E����of��A�[�f=���r��lw��{���Q�4���戎u���3u�LT5�-��ж��0����K�u�e��yʢ�m�����L�%pb���w�lƏo81W(6�DJ��s���m�`����1������[l��y��juˋ�M�0�G:ܻk�L�*�c�D�钛s�ۓt��¹�0�\a���|)�G�ٗs��s�ڳs;e6��6�m�ԵV8㜕A2Ŷ�32��r��p4lQ��ո8�l�v���V[�\eXʭZ�]2�.L���uۘ謪�ݺ�q�*\��%6�P���[��fCS���F0[�.���\U�U����9�4�M�gc�.(e�L�Z�ԹD�M���3�c�������1bڳ\L̦n,m˘�UEe�̾�nY�{ܴڊm��S��7.�\˘�����Ɉ�q,��$���Q��{�.�Uv����EkoeĦ-.m0��幎۔�V�j[K�feiU�����R����nn��\�;{u05&�]�yͷ70�QS��e����1]bvc���j�lZ��S-6�j�A;��q�k5�K]�7EL�c��;�u��vuwʡ㈯�u�£Ւ��<�\�b��A��q\�1�U�������R $D�P%!E�D���u�}??I�t_s��=tS���|�}��������(#������~W�}�����{���������������8������� �  K�_�����=�N�ͳ����W�چ�A���ڣ�
�6DZ�i�+)zY����+�����U	�[�o=�5���clw�{!��y��J��&�k�NH�H�A�7� �x��aC�]]�@�n3�|�{�u3>c)�is.U��R�TE�i{���D����罕�͹|�������{zq�p;�޾>��SDY,̃P�h<rڎ���[�(Y�C��fͅ��h�ƔQ�T�xn������B�vO"V��	5�/+{Z�0��W�z5��s�M��ї�����I�-�����M&!M���UY�^�����~)E�����Πk�A���.�#ڵ�ψ�LUc���h>�$����zh�	%fU�*Z@�s��!MH���K���l%����b�4�/.n�qzb.���Tacֵ��g���C|�mU�Ez��D���ֲT.��x����v���1d�)���1�$̅�zf�N�IBs�zy
?���@S�nZ>h��Ö�o|]9~���I��8����I��z3�>}x��'(^̘1@L<�b(�����F �Rg�i�2.�
�\IW�p��%^q�ՠ����V�'��]B��t�YR�n�����A$q���k^��"���r��b����H���P��+15͞R�}-�;��"�&�8�c��( ѥzg&�n�cѪ7��H��e����]���V}y�tU������z�N�{\
�r�������rG���۹�	�0j�(�u�V�E'9�NW�Q#��ij�
����CP�7��G���P�%�����1����	����ׂ��k9�׉��@���X �����b��nni)��N]���wY�J��	�鬤�N�Ȱ 3�#eЯ8%b�H�����Y�zJ��<w��n0�%ݷa~E#�<� nr8��s�ؾ5N//Akf5쉄�q�j��%�{i�[bhh�uS7�frO�G7B |R�2N-[���%��?.�H38�rj����c�$6/��<5!J�ӊ|�Shx�0N0���`X��2ku�I0%����3����` �݁iQhT�y(2񖒳\_��ǯYb�#��   << �  ��t������������S�l�E$��I)$/�d�)�?����("�BIH���e�|g��v]=����'�v4��{3!�����)�?���<P�[�`�r��ob��m�����ڥ����P�!�/�9���@q�_/�|�Ed�D	��m��M��E�
�̛%7�w��?�/�[��I~�A5%-S�4\ђK	��O�!E�I�SS��J��6��y��x��~�ǳg�m ~q�&�k"g*�c�R��ST�ӈ}+�^:�QLe-7%�p���7EeáŎd)���8�JF��?Z�	3�0�p]�$�������k$㜩.7��NwvA%#ZE�Q8GU�Bh�[�/^:,��5�u�]D&�u-t1N�^3t��C>-�S�$5�F�鹡g4�H�BXE$��"�]o,���� |I�xL�QR_j�>%4�<�R��U��~E��F:am��`6��5iZҺQV��VI�F���]6���x��]���4�"��L�����Z���H�6�涰e3U(r�CJN�"�"K�{�Q9.�@����Q1�dd�	\@����{�x�z��,Z%W	����aN�1n�!+A H�	A���F¤fn�^��^]d�h�����i�D��,�L-�ѷ����N���<J*��ba�P0��=����,�
����i�����a�(41U�YP>��	�Fl���KY(�4��@�o\��c,��ɽi��l�Z��M����KAC\����}.��M�.����>a�ی ����ֺ2̼��#x��CSA���1n�`F$�(�x��U�V8('�z&F]ʃ��Y�Y�6@V�c͐v͸y�\w�-N)[��9�����]�>Y���E�<#�F�z��n\�_��;F� �J|��&�_f���4�h$�	�ZR���ܻIO�iG#���E9-A�"�LF��,S
�!�r^�T�`���.�b:��*k��$���du�B"׌]$30� �����b� P>�p��pe�b�廴���J�P�J���!Ѱ���b�:s�Q��E����� �|��ﱳT藼�/^&�ǭ�N�t�tb�ee��6cl9A��a�[�>Rm��nZ�&�.��s��Nj�+��XF�a�! C�9�IN��C�.��0�.d"��T4��[�����"�XGGd���?!K��!}֫�2�c<��*g�_��i5̵Z� ��� "�&$WMu�S��sT�5R٭N�W2̢�f5��f�l�6s�ʺ:�95m}�ۊ�X�����ʻ1;��~#�!�jθ��3jq��T�Д@�
�OP� �Na�i�u�YPq���=?��U�99}r�ꝟMWԆ�Tw�bda4�v=�28xUoQq<��y��v��H��,�)����d�������*��c?~���@ؘ�_�r ��C=u ā-/��� O�s�.�f-�w'�uN��w��i��ŽI{�C�v���9�^����f�8�sg���x�`����w�/N��|.�^��'�u��eq���:�yy�1!����%��R��xz|y��X�墇Y��T���Pz�һ[e��mV�;�6e��)��sې%��" T@FD�U!	��`�`I"8�E%b�El�ݺ�<�^J����?(���Q��{h���X9��W��w/*��/O��������evc�\Ֆ��=�� )�i��RJ�
�nᳫ���lo'#���;oo��Uw�;^^f˻N֤�Qܪ�C�fy3�K��H�G"��G���#�C�u�up���{�b{��Tz �Ҳ�Iz(��;���=�=X�6�h|n�����wb���z���U��Ǉ;j�]h�&��)Zi�-��9�'G~v����:�*g1f��Z	I �q�LaR��/�*�B@�.ڣ$R2f\���4#����["��Z�9<:�tֳV�m-����(��^4vI 1-�$*5����s���o��˾6���T�y:�ɵ�ԩ�Sa��- z��`T	 ����䟄�z�IBHF)!�
0F -ae�UAY9��s�nt��Y�2ڧ�Y!	Z��"b��¦!c�9$��Y�3&�$!�_���$���I�vVI�QX0gm%ƪ�fn�s��W1�b�#�sR�� a�+		�Q� �BԤ*
��Ls6��5̔8�5FcDSRQYr� �I�-�z�լ���Vb5�̒�� ���
ȘRIEF3p��>�p�Hc$��ϫўd��d������HH��ÝЉO$�5�� \��:I�U��T�R4�4;u��Ur�cQ���&qr8��r��3������xi�a�V9QU)�G�ʑ�D�Tl��l�D��4����٥	UU�B�J//�I�RC�*)'E��gѦ��4<�E���٦����]���Sw�e�{��Z��2��� �j��2��\�H��H��$�Cß_>ZgS]i��2�]�@��U��K�$�1$���z�L�b�NdNڕ;�Tؗ4Uv�U]�K�Dxj���.섧4���5�ʤj�.b��A2$\�P��Uxb�l��j'v�9� ��*�c�f�%r�����Ma�[TY��C��P9�ȡ
�P�1�X���g;��iiD�U�c����u/��W�:��;h��A�3�j��M}��7*wU�hƶ�b\���M�s�*e;7+��7<��-z�5����v��-�2۶�ۻ���E�Kly7
��r��w9��8���^{�Y�o��SĪu��;��ίcD�)[R���k��5����Ysp֍����u�nZY�qDT岽��v���Q�W�9s/R�aN���n�v�L˯�q���,f۶�����p���w��և��<곦m�iO\9�a��W1�}�M���b����o���}a}B�[��V���{uث����^���x\2��2���
�X.�S֕3���Z�2fbU澷�[�c�'#�pĘ�d��S����B�V�z��e���0O\�MR���6��W�,÷M��e�q\���Ո��6댻�����fS�8[B�}i��f�fg��ۡ�n,Z�_o\�l�Դ�^jk7s2�H��7r�*��mR�1*v_u���꽛׶��(�\'4[����*�mk��*�n�g\5�L�s�x�cZ̗ƥ���Gn۝놊��Φ�jk�v�.ړ���\g��i���k��e+K��C��f�Դ���#�]�-�f\7��ε�����of�j���JmJx��@R�}ٓm���q��f^}���i�
��3mM�T\��.0�a�#|�����}�nJ:�\onG(�U�}�k�r��4Q}k�ݺ��6�V�{|���eu7-��;�}��|�3�/��y(��nDMe]n*[AR��EƗ0�Z��÷2�{ٌ���γVs���m�M�Pμe|��-����M�M���n�t��&�v�������ƶ��+�ܺgi�Vڕ(�t���;�q�r����uÄ��r�`���q(��c�C<�v/
jum�����ͷs���D�B���g��Q������q��\J�iہ�UnW0�1�\�Am^g�b뉬��6����g��m�ٖ���S�2�<�dF��nڕ�e�\�.0��d�wo�)�s٘��&���Fۖv�5=�S�2��-��w��������-3͉�Fو���K��y��=LB��hs�5�/F�/���_f�%<��<�0�\��fgd�s�t��n�c��0p�M�I����(�c�.>K�������Ά��`�%�c���Lb��19*T�mSל�֪���႙Wp�=��_W�p̥tK�+����P��Umv��t�
�=������y�Ɏ�5�n+^̶�(V������R9O<m���^��F֨�վ�����:��ge�)�����\λ�;��{�����d�b0�0�-��v�-����q�ȷ,P�151�}��<�拖h��;�]p]}�:�P��8�\[�Ͷ����/m�m9�����r��oos}���g��AN0h��>M��}}�UK��]L�ɉ�}�մ�;�n�n3�Y��tͷn���m�eSh[L�Ɣ�*V׽��L�䢅����\[��n8�l�W۞����BڝpQ�MK�-�ɚ�6�LT�q2�������ֳP�+hw�<n�$�Y%O2��$Z�[c!� �&"�(
E UCR+ Ĭ!X$RVE1�Ʋ����G,���d�ԁ���|a7�ɨh�FAa��	��Ԑ�� �C�O1C_5�X��BgU�%F�+j�Ę�ȡ!Y�{l&[7,j�-"4����T���G��{YF�Z�f���kV�636&�f�P���@�)P��b)b"1�*$*[D�()PT��,r��f39��g*��6�"�H��C��j�����"�,�H�H�TVJPQD�EU`�UED+cb�EPQ`�c"1""��EAQH�b�,APAU�
����U`���"�2�)�=�����sW�$���^����:֗��2���:>��w���������y�������uo}��w:�S�ф�!RB~�dI&�$��t�{�B�x�q��_�������(�Lr�s퉛pDQ?9*��1fߋ5J�Q5?�W�o�1q��ÐH:�\��)
O�׽�c��}���?�?����>P�?�PP���[}<��m��6�mHm�SeG1sl���G5B��1�\�sM�m9��Q[IK�%rm�s��mU�kfٙ��[Vյ�6�ʲ�-��h\ҙ�͚lm[6[�
��m�h�Ylm$�S��؎a̩@,�� ��$%�I��/�EAE���ADb(� (����"ň�~�f*V�cm�p���Un��C�f�֗YŊ�)�4Zb�
kf���ecdL'�	�$*R5 �Z�-��d������R)IJ�Ql�+`�A�LU�A(��
��Udbj��l�mݐ��L�С*b)1��Ⱥ�RUq)l�5*�F",Q�6��X�(���X�U`��̢:�E�����PA�J�$\�.ci6���{YT�H�`��Z�VMjE�,����mH�E�(���:�DQF�QfZ � ��c��*(�B�+`,���*��]묝�u]��\�&Z��,e�/��(�j�Z�X����5��dEH�dX�bAE
µ�*�&!RCP�!�+	2@6(b��X��v��*�q�,��UZ����2Ҫ���X�4QIU�d��	 H�H��+��~>���_#���?m�D���-�y|��w�,���w�q�r����y�^ܱ�+���~�!��o�T5>q�sټn��d/��[��������tN�F���b"���iݨ9�t�T�]aֹ�ȱ`s�T֪+"&�L���H[R1R�EAE�,b�1��}@C��RG6c�8� ̯���4�.q�����+��kw
��4��~�}�,|��o�����!1�ko�"}�O���S��&�|�x�z��{O.!Y�].w[�39,����E�	$A�$QM�*Č���QI#����R9eW��(�X��Yl�PDU�`��@v�d�%`���9��\gm9�6)�hL����M2�E�;J��n�X�h�A8�(�ER �m*��PQE+A	-"�������&sMsf��&��װ�2Y�[e�4��F9���)��赀v�Cə�2'�X$�N��sx8YI�/7)r�i�����_��VN�{t�<{��9äQ_[S�*S��}����0��a�|���Z�x�K���b$!<'l嗊��Z>�W�����T��$�0��1̝U�X�����t�&�1�;��Lt�;&�l} i�0w`��/�&�'��ͺ������ޓ��F��F�
=���F�q�[�i{�d5��2���B�7n2���<�����3��)���<�R��+�7�>�^�cr&�T�w	�w�Gq����.ܝ�B�R�9�\�KM�`���Mw[�W1- jJ��������#���v�BI�Rcg,��ڈ*�T���;�v��.�*�"�jp���`yk�ްp^[8�x���D�J�O��<��`�{f6��,4��Ý�B�����;g���wL��h���BH%�ꁉ0���4\�'���C	���"Z�@���*�e>��8:��[3����86�ݬ��ÏIr8t�U��i60�ߥ
I�%�KI�4���Ξ�A�Zk�@hi�U�Õ9d���c��3K�98d�P�,&�@&�%���-@`]Z�aM͆�&J��'G����'��>�wcL���c�̭$n�ֽ��.�w�Nb���`d�O�p���ߦGY�{�)��|�s\�$��J�遖4��o�D,�M��wT�fN�#��DdF���߰UݵrIYd�	��{V"ռmZߘnt�0��8�4o��9��<�mk�bgo�.@����QR�T�5�6�(oΧ�����6���JUK5}n�P�\ѭ�m�˲GJpG w�Ӳ; ��K�}.��h����Ew�nܝٲ��K��r�s����	=��ĺo�n���h�)�����{��tn+�R���$���/���"o���:�ɮN�␂5A�l�y�_v���OW��Ld����r��\�k���;�X*��GU�]�ը�U o_�p�ڣmE=��=�z�8H2��Ѓ& <���l��/����!��]i��&`͵�ł��V�L�"�A��j "e��,Qb�°�"Ȣ�,�^��$�1_K�ʝi�;IGpw���Ĩ宵���U����DDTc�D�PV
�V1"�Jh��c	��MIAE���RT�4I@,
�J�[E�Ȋ(�"�F	���۹�X����]���2XASF�mә-�i6]��P��� DX�U�",-��[�~Zm�EG�,QH� �|��rBV*�Y �H(D�a�:��AAVbjdMj����V+YYU$R+l+"�`
CP5BpM'cdEE�sUR����Q�U5�Db��%E��5%�p_����]�{)*��/f{�S���nֹ2k��Bl���}������c'��?�V
ڟ�CQ[`k'bV�2W��w���9I���[o/�>��x9_��ZG�Зw�c���L�?
�9�u���u��������%�QJ��E�.�t!����AR��)���Hl�e&��?����_�5��O���w�
��ݹ?��?4*���Na?��E�Mm̤>2�0;y�F���6�j���#8;i��
(1`F��g��H�S����ef�u��$\
T��������=��MC��&p�>��c�&���S���lm��SY3��_U��L�`�*���ꉡ&�ᜃ���e�Ayc�j�p`[��'͢�����M�p��$/)��)����`ͻFsbϷ�@�,�*�P?-Ԑee
(Œ �&D�)��i�ѥ$G "�/�J��y)����"뚟+�g{������V�J�8&�<35��AWB�l��*�B��PoH�Xl~&����l$�Q"y$�d#]�5D�%�s�{����LP�Y,JR>�q����y�xX�-��X,�F�|���¼8���i�v�I�Xq�'h$J*lw$G!����G� EAbT ��1FA"I��yN��/NMM��8C�D�SC2;JBb�D��vOiߗ��wz|U��+aǾ♾�ǽ:�!�p[8(h4���(���H8@���L��[�݈�r�m�9��,A2�:�j+
,�)s���f)�  yu�[M�l�bG����*'��@��?c�m�PE��EQDAH�V


�Q��QH�d\jB9d�cLC��TA��h�h�w\q������A(��� �P"���%d����@M�,KyȪ��O[j�����w!�h��!+7�%d����[e��N�����1T��)P���*¢�$��V�X��*"���UPTJ���,�"#���?��!�'0$��PdT`�U�b��V �6��Z�6�7,�X����T#DY�E��*H����VE�KaG�d1��Mm�Yaj*ŀ���]�`�� �, ��J$����aé�z�s*#I8����*�=CX�,�aRӳ$Xbc9�z��ÐG��A@��&�O��||���,-��Z6�QE����В\?�����i`��ʈ��UYQB�,dF(�#
(
�PQ-%IYKT�
�Tb�*�UU*6��26±aQB#��(���[`%h���.L�0P�6U�TK-J��J@m�	Z�*�DK
��mKKcI%)D�<��C�w��|���*���=�V�~L
��æ%����/�r�1��/����/����O.�N�<q6mx��Kn�FXUe�F��H�B�������	P������)0�O1&�&J�X��c��T�v��}����IF��,��F��?a���z�!b@�e��+�����VM��,�%N��vt��b26Р�5Ķ���AR%�~�þ[ ~����:|�s�]����1bL�b�Oݥ�M����eй� ~c/��?C4R��9� B�Y��d���n�:</2�Sa٬;��/�9��0�K-�(|���	]f�e1�ֆ5u�\4��lU���y���euL������K��hm���,A%��W��� �M>kW)N. �X굾���د�40EAߩR�`��	�XP(�  �Q�UJ+(�X�b�T��mm��V�R�����31����9caթ�Gskg��4v�MJ$X�@X
�S-%��B�v�V, �,����"�XB=qR,QAEER(���)$��ꊹ�6�cjm6��6]�W~u��m�`ٵk-���Y�Ud1* ��P&!X��T�
� )AB�b�Aa�*��g[��X�"1q V�fXJ�!I�¢�P�%J�(*ɨa#h��`I�QUE�EQPUV
�R�AE"�FL�[��.���;�9���9�ɚ�6���[L��
HT��5UR*�O[-��)QA`�U �X�)1 |�@�т1dU��(��D�(E�s"��I� .�^�E���"�ԕ���[J1d��()9 ��E���]J�*�2�FҺ��&��ڭ�v���CY�(	H�HF#�Z�"�"��T�s%H
��%I	���7A�,P�YY*�:����c#�a5�Xk�Ke�&ҝ�sr]\�u�m�PR#
ピ���UA��B*Hc"�P$ a,*������"��k1(�[iV()��U�:��
u�wj��f+j��QW��X��ٹTcF
"0��X]9����U;�u��W46 ��id��2�S���-�����$AUb�ȥI5�!$�C<��%HhNH��W�c�
��X���[�&�w�A`��U�X*��V |LC�CP|d��!�M�P+'$�Uf[�ȌP-(�FE,��cUV$Y�C�J� �J�E�I�0�
TĬE���*��YQT�V��3m��Wl\���`w��6Ts��.�;ke��-�F,��AVVJ������a�(�QAEA�Q���j(b�1!}HT��$ o�'�
�`�I�q"3YX�����f�` �.Z�Q�X*"cA`�
e��Nm��4�*v�9�G%ʳ��*LdX,�`�0dQ��M��D���1V[b�PQAQQT����KU �����<��dsR����w��s]s��7��X�S���ʋ Xł�X֋"(��YfҎ��"DQDTQQF��$R�d'$��NM@�� �"I�E'�H�����HV"���eE�Jʍ����U�AU}�%�������R����'��?���E]����N��k�I��1���Fi��zj9��0�sW0���a�h�Y?��AC	�)����%X��[X�lA�1D�UX�,D��YKD�QDUE�*��-�P��Q�*�F @�p3�/K�P�5}L�{���W���n']��W��5~�q����_s��{Oq�l�~o[�m�ƫ����7��=a�	7M^տ��kնݧ�U�����x8S!)�~���[]���X�;��IT��/��ߪ~���	��)��o�5��O��	m(T��?q�߹m�q���	Z|��$��|�ŤX�{����4��A��v�'N��4���<l=yVA��W��^������ܬ9;L:�/����C/Ά��A*�����l����;d5)V��g^p��J��,�cc���_gßEQ��lj��?S��p�k���%՛��a��s6�c��ϰ��V�޹���U���Tk�m�-�;���y#z/+u"J�fR��x�}(Ǡ�^E=��ݻ���4�CAA)7���w�`����	�Kw�P����f� �氥���N�:Δ���5�qx�4 Pi�%C~�p�&D{�M�C��/�獒�U"��<��߃�uKݧG��1���`w��]��e�H^�D���ڣ�h3f���̸�=�P��.Q��f��.���/�>�! ƚjP�9Lh�C�8��cQcL�_��*�����h���v=�����M���Zf��X}^{��V�8����p��3�������с�O�����^ںɜ��9�4vY�s�����R�}A�ҫ��w�` �O������1���r���Ⱦ���iM��?7��[������S��&�8��R޹[�{6���8Q�'�a�L�@� xxc'$!)�ϴ��[�px���[u�3�xEP�m�ጺ�]�n�<��~�����`�BT�I��F} w��z�ȶAҨ>�ԝ�j/f��.@Ɯ�gw��I.�c̟ǃ	 R;�%ϱ�3�C�>�	�驛���D���gܾ�r���G��%ڊ��RM���L��u�{�<P&�i*���gq��1s1�!�;�kC��V�,�������<��c;\���#�VJ���\)aз����̵u�cqV��qnl��&D3/Lx 3��G��aS��o����t�;=���V����Ǖ|���&�|D��ǘ�K�J<9=�Vt�3�M4�P�s�q���E�ՙ]�rgx����I���'����A�K�*�|�֙�>�FK�$%\%�t�Ҧ�	�#ϵ��Gy�q�.��vQ6��)+7�]5�=�͎��VK��Zq�u�nT��N@p�w:,˨D�8�)�0���ʀS��)$�$�����<QZ�z8�K6�mu��7k�i���ۭ�L�ߞ�v�u�6�wg<�1�Y4��	u�[�˖v��q)D���n�~�U+=�OrF�V�9Ɖ�w�HaFBv��.���>�"�Ŗ,�5�,����cJ�,'�An§�?$p��&u'���DJ�n(;_�.� �N�]�!���ՓƩ߃w.����� �9݌H%��k ^gr�4�%�dIu�P��v=��S^�J�Y;1	�_R �	����UtK\q��@[��9\��=���w#tx���@�쁘޼������!DgG�>��3�U.8$^�j�Gr�͵���B�fon��Q�)7�W���tn�?9�iv^���E���d��������h;�Ͻ�q9�����6�������hP��6�q��Էj+�R�$�Γ�)y�c�<�8ۨ������-�.�:	!�ܱ�[ѡ�uⶊ٪�fN���I�a���E�1^�J�&��H�)�e����|o�4�͙���ze��Y|��t�<�CwC5�ZT?iKQ�s��G�gvЄ�^��,��M=�AUP-=������ON��q���#��5r��쎓���O�H�<�ڻ{���]�w,�U������&	���#�kO�MP�_�&��1#p�������b�`�E����o��������R���pmjri�w��)���&E2����2�}���?����~�w|UӾچ8���I�&�)��p@�@!ٚy'mB���TV�����D��/�Ƃ�+��L�-L���:�x7�%x�4>��h�H�e=:�O����7�k�_������g��iLH+M��<}�E0D�D���0	(^�,%��@O�'�&���~�s��-�R�"���+p�j�ŰV�NJ��DM�f�j8�f�E��[[��\����삻����@�xȵxH���0"� ㋶���Щ@y�v݇�V�gx��	��< �)��,�A�i_׾�[�_�?6ܱ�����S�[��.�Q'5tw�J�MC_<�φ>��M��.p�\_�h\􁹝�TT
5��}G�F���P��IU.q��T:�B��2d�`A��dA�'K@�pH�;��&���%���&��D{	�f�eS�f��N�����\L�x��p��׃u�w�Ӕ3�㺗�x\��%E����Y�Z��;����=B&dN���m�ٖ68YHE�C�p��' �j�P�ٝzͤ�����}u�@�I�݃5�ֵ�3��5|]j��U����?'�i���f񈖔���C���E�G+��j���R)�(b
�c���+�mE�F8� *��#1!X�X(�2�P�3Y�]���ՋD�Jc�%�d[�K��ƨ���(�0�e�E\�he��kh�E��ʢ6ؖ��Y[Z�X���8`婔��l�W2�m�PUA�
��ƅ�����=0X��*X�B) �"�"�Y��`�dd*�DA�"EX���1b��b�T"��b*�b��(���Pb�V*�
H��A����(��F"�E� z$V	AQ�fm�f���m��[%E�, ���Q�����*$X�"��E�EDX,@��jl�mLͪض��lU�lٴl�6��ٵ��"�RV1c 0"H=U,����&�3g���ʻ�w+�}����{Q��1���/����!`��BG�!��P�����d"��� *O�D���'��JF�
��v�%�M�i���Q�����~n���A"V�����H��2�6ڣ��G���Dr-<p&qǁ@���_2��xB
=��(��	�?�P`�M�V� ��
��{�� ��ω���=�}"�4�+?�+T;zZ�mc<�U�9�R�?� �l�<�����y���A "E������A��䜹�d��CS]UUY]UTUL��v��ۅ�v�w�O���H�W��D`� ?5"��Z
E��m��5y�_�����3�9�sI�S���ck{9q�l�M���YH�$AT�U����$`I	2,����s����鴟���r����t_�w�w��O�f��{Z޷�KM���o���>����-������|����5څR;Đ��N���m�t��%r�W-�2��H�c�a����f��i%��ҧ29����s%6��#�eQ�@�Jm6���5NeK�W4�jګa.j�B���-�أe-�l7�B'E���15M5Z��Ϗ�?��7�?4����	����#~���~G�/�����?#��z�XJ���і?ܧ����xx%�~�u��_���E�Z��It?�{��v�+Jz���[)��?L=S77���R�E��8�_&���|z���O�t���+��S�s�P�ף�� h@�� �s���M�?]�%N�_FlM'�s�Z$[�j�M5�6EF��R$ݚ��Zd-w���Ĺ\�sOgR[�s^�<�f[R��'��9���3��jOy�yf�r���_�,¡��H*_.JčA�5�#�`��/�c��DU�%a����k�Q�5ËG
��<|�16�=���xD��"z$[��GD�����?H��"z��M��hX�/Y���E0tIU\٣E�`��ٜ��^Y�Wd��j>b�A��t��D����۸���~<V���3����(B�Ƈw2+a@�1&p�;<6kFH��{�i�L�	� ����U���ZF�?��;Ω�����~�
3U�{D�#��\��S�YF��u�>|/۫<���1jW�|C���)t���)����m��,뗶�X]��eS��z�"]�t����p�x s}!�u"�;��}�����kj�s�{�F@ܳ_������sYіʨvz�R�z>zl��p�3p�4�\t{���	����͵'gR���Fv�^�8ىyeɲ������Vl�t�"�Ÿ���R������V���ŸV�-��ሁ�aϹ�JF�Ǡdۇxp���wF��D�a\�)ϰqt�#ٮ�5��ᄉ⢸�(f���݀��M<9�c��ii§jn�A���4�i����P����hf2˧7o�-A���j=ZĜ
�DY�|���v�߹g�>4\h�c�]�lG���Gy]��Rv��8��Y��P��T3q�*�),Yp��A9�|
S��%LLu=��K��B�l���	F;V�4��I�X���Y��I sI�9�UGR�3;��}9�~L"|�.\��VG}���m�v��S��r����ؒgf�&	6~��K�v솲�{.��*w�+���xڑ��x�#�8!��L���퓂 x�⋿��'I�[��׼@(�����[P&�m+[mk�w&k�H����w��Z<ϻ��:dA�t�QE�6��:D.NdVp58^s�D/���H��Kٚr���_= �z�oڔnَ�hsf(jn�{;>Ϣn�14M8�ሢ0���0� � x����Y�d�U^we��t�C'z���F�m�ʶL��x�A�/������cR�!)#�~G�`	k��:�r.����5���+��i~i���.��7.�j��N���>��݌���v�F虑���K�}��in��)�B��O��S#�����gv�k�;��~��9����Y�����'V����	�]��[}J*��VX��Ռ�&9JO�;��=��Y:('���u�J�3�s��&V�~9�H��p.�"U��qr���
���@s��$��Y@uFxF6aQ�Ø8b�bE�6"���^���ۗ-�׼����׀(}Ϊ�`J7H�>��I�d�<C�`�t� �ED$Ȯ��n�.��#H������ԣ)RF#4GMp.	B�[&Wp��,�89R����<&��\�����[�!�㢽0[=ӡ�s~�ݺ�]�Ot9�n!M�&R]�ޚ�&�BJ]�yb��ڪ���H��̀�HZb�N�b���ϛm�R�0�.l������Lǧ./�yq��E|/�6J>�ѥ*���TR�׺�n�rX������:�A5Y�9��m;ԥ�B��;w�c�?X�'�U߯���xsN�=�yj� �G�oQ  � "���!��~��gꟲN��X���R|�����m��M4Ak�6|���m-m�3i���6�!!�$�a�E��x����w[��w�����\�W��=���쾞�����?�yk�Ϩe�jI����S=QLB��I+¦J!¡�L���20	b���{����x?��\������+�X�����./'VO�ק������rvbr�|�-��m�r�g��*�a����%ς�?Xݫ�|��&fX��Xd�;�����=$���_f�y}��]�C�e�~V��	��v8}�?���QH%�	���$+��?q�����ǧ;��&�R �H�[ز��K�d3;kEfsK����3��%��_d>�^�!G!������*�]iZ�2zrR�>�藎���l^("�� ��:r��74��귍ң�-���gH�>o��u6�F_8�2yI�j=���T�<l���u�	㪾��B���Ӕ��0���:3���1���ω�!�*������l�:~�7.�˲�9��!04.!��Jq���T�95�ɺiq��R('D��z�Wǰ�C(�����R��$꓂�!e
!������"<*�Y�t�* �V��i���M���p9����mgt��$��{X]V8���:��,{�2���rg�ݕn�y�Gm{r��O���I���t�P���GF��7��E��.����`D����^��L���>�[<��'M��#Nօ���	�Y��d(�3�bq����߆;d����a���;s5-,婜����x�6� ��&�8��,�K��vHG�ň�!m�Sd'�ټ橒Z�%3�@�ukk��A�,�lj@UR��J�ӛ1iր��|q� ��A��� ��G繦yvQ{R��Ib���lٮR&����Gὖ:��WjH\9��Εqm�z�l���s{��i2R�s�Vŋ����7I`�p��$�
.���8��ʸ��Kę���/����Z�ݎ���釗���g���b�����j��7�V�3������Uܻ�"��u%]��؂Q��ʪk��H1��S�&P�H��G��'V�*OQ0m�w3 �$���KoW}W�,8��	�D��vA�Uцη�
�h�˖�МnLK,�	v��-5b
���Kėx�W�}(h�J�(���=2km�"K�hN-:���?<�;���)�8�-�K���@4p�z�Ed�X#�Bׁ� �U+�^\�N�D]��p��l��*��~�=s�c!�b�ѡa�,j�v>uk�6���9=�m�,o.Tl� �I�ߛ=h��12&6�&Dc�t�g�s�	�I�&,r�E��j߹���`�m��00�|��G��aiuM��adAv���0������=�������_k�H;P�'3VUŧ�{�$��+{��E9�-��ǅ
��?��-s�{���X&�-���3��cE�%�8of*�g?�����-����&��&���~vf[~��B�i~y���p�=��~	�����ۋ���^r|oB9#K~x(1o���ы���t�I�P7�2*����{k٦�PgI���= �����O������2/�$�vf�I���B��4����A�]R�U�^�
�7��(dz�,�7���hNz})�v�b�M����r��<��%���7oR������B��hPC}.,f�]V��4p�3�z}��x���|��oV���^��ݽ �%���������S�TB�[��ֳ��)r{��6cl�Zz��C�OH>p�:��l�E�5��3�EJZ8�*�}�k��H�R�PN�{���c�:�z��b"�(ǘ]3OHW^
�1j��*h���vH��CMW�"����9��d5j�(
P
�t�Pa եOe��m�f�ٶ��$�!"B%�n�����G����+��wnO��8�_�������S|�����WVP�Y�YQU-T�� n%�q;�{9]Vo���9B@��'������g�ݻ�`��<�x�����"��>�5��_� T�������� #�RB�#����?��<�[v�\���{3c#o�ޛ����f�w��	�|V&�N-|j��N]�+���#rXke^�g6�	��t���O�Nq�  �[�{@0�1b��ҮI���"(�eǘ�<@�b��}z���Á�腊L��g��b�!WniD4��o�`�K �c�.dD��Ӽq����vm���|��f�2?s��0��R`M���:cV���m/:id��.�`a��X�qg#ˑ�s�94A��pK�{O�fB���������
��%QE�C=�#��3O^���F��i?~r?ӈ��<�J�6%3�vC���[�K��}Y�6�ܗ��}��u s�b�V0go��I�G$���]��;�	L5L[�EÀ�C�aA��;�0�nG��2�j��G9COT��)�u"�8I�l�-�E��'ۭ1��,DxT�=�^>H�� חt��4]��yo�|��{�����on�O����N)`��e�B��>+�y�gzf�.KLձ)o��ѪrR(/|��7��4��*���^�O^Ӕ��'�A�Wc�-�BCF����;����N�$N�~��F ̥�iλn�vL\XX�q`E�&oqΑ��Ҋg/�(\/&��-��uN'u����R7_��q:�(��]A�`o��AI�f�u_؞B����ݚ���q3�|Z#["���.Q�hM. ���BN�a�i�e�Z�4h�E`>HD���=�z��ol�����a�6Fp=�֧$�`u�I��p�J�@����Ȅ��8��1wEԽR��Z�ɮ��o��<�d6�7&�i^�^T�{�v���9�>�dbKު����q:vYqa�X�������H �V���Ϣ,C*�����N����n8QL�7� �S�8I;��!�ĕN:a�q��gr�e���d���[p�Bn�c���;��pl�FMVa&0����Ny��v�˗>����+R�n&?&����~�d���L�� 5�H>t�z�]rW�gu.S��0���Z��%u!$��������k1K���ڕ���$�-�W<��=A<f�
�1B��OB�K��	-��æM�����a�˘��4^�E��5� ~�8�V�F����pZ��@.�F�[��&�)!ƈEO�-����`z%�I�'s���9#�r�69�t�u�5U�����L<���&�x�   x}w��j�<h�!�@�T^�|f}���p��A�}�yD����	z�G�<��U-�����*�RsZ��(D m2�_��C��[�*1�7|XZq�ߕ���/R�+����ڶ�]V�`�ҝm��?]�-�^|�����?}���Ke�{$��b�h7�]zY���E��k���=M�pM�.J����|h���7��4�n��بxS��f��~y�r�'�4~�N��F�z��V6%��	�{��j��Gǯm9x��17���W����^뇦�o��`�����I���h��Y|PV�8xxRr�
рKU� ���-�)�86j�-�ʲ3uBJ]j�8tC��ٗ*�r���
?�qт-1R�O�)LCh�o�Awb�Rg�a;5R� �>�ª-�y[�y���:��o�����7I�A����fo+,�6r[[����gd0n�y4l�ҷ5�i��A�H0JYHb�>��iZE�iK�S:�#�u_.CY>^1�l�}k�[��s�}쒗�{Γ��O˾�~�m�m��w,i�"�6i���`���͞��5[mf6Y�hDu��ٱ'��~
�����N��v_s���,w��>f���<������9^�䵔�_��韀�[�bW�����Lm�D~�����8��̥�����79	n�*��im��*:S��/��~Z��
������[����5`ַ{��b�[�}wk�_�)��=������(��!����Mgi�n�v���"�Wq�*��FDCٜ���M����ż�j�r����!��\u�X���ȋ$q��S��/�I8L�Ȩ���*p]���Cm����#/khh�Yڠ��ۃ�:��!>	_Rޚ��(�S�4d�ڜ��^���È��F��31�bhi��U
1��?)����m|��WK���ȏ��W�e�{���
\�R����U��࣫�����cp���_ց�I��� � x�{�{Ϭ���׉��~���7��>�ߥ�@����ܖ�]���g����b��?m������N:I>��2�b�����&���������O�`�aL�{<���:����}��2?@Uc)�9݁�y��>�ѝ�邱e�Mv�I��S^�u�u��b�!<���(���ϥ��T^sL�<�bO�ɑ7�bZ-�>((��sv��q��q�6{Ш�lN<�)N��/bc�~k�x���q�A����:�3��]��S�DRhmm���/�8Fk��R���?*�Ŗc#&��pa��L��r�G^��41��۪ψ<X��58��E�����1Usk!u�q�{�o�4b~�9�g7f�=�'r��x�_�4)�'��r�:j��GD���a)l^d �Y/!1��4fb�1qw>��Q!Y�%�Զ�Bn�C_F�HLn����ѦT�%Q������hl����ؐMۤH?x��֙��eF�0�sѝ�O�rDLc���!�ó�-��k���}r�<%��*H�9\�wV�#nq؞��7H0�Ҵc62�b��[�J�*���hy��zٯ�yߥ��S,,� !�M����=G=���l���<5B{�w�Rݜ<���h����PZ<�!�HY�^��
�C����Cx;P��,���9��48?T.ӕ�ɗUvTm��:J�x_+3��,��8L#!��#���9Xt$-e�|������3c�{it�s�"����3��@���X�u��sF���C0��S�g1!s�$�b��ʓ�bmM缥�y�$����۵��8��Iᨆ�E�j�Gv��p�Ԇ)���_����M�<�.�5��	�~���8�,]^�.���H����c[:[b�#.6���ojZ����o���Oa0g7�������?p��޷e������V�-͚s�Nk�y�(!ǀ�m�x+ܡ# ����eO_��a��(˽��א�k\[�,��$�����[�W&q�}���xj���۪��4t�:l�>�Q�r�M��Kͼ�l�)M���{NR�����5��f��ݺ�:��>�a2e_�c��VM}8+vr�W��ӓ��A��%H�d�h�R����;3��M�g�nFwۗj\f	;:ϐ
���S!>�;��i��^���kL��>���Ow����(����C�8��s���� �=ǫ�K{���d�b�"��s�}��e���Q46k\����wNC�����r<K6�2˅�=�U�w]�k8XvbbY���N���EPH@�4]( =�����֍_��S{p��7O�kk{�cO�a�c��X��ߖi�c����r�����Rs�^�`(�o�!CI�s���2盪��`�s4u��+�T�ފ��9٢m�8�,m��JM�1t��EAPSo�6������nQ=jL9�m�8�ߞ&�ϖ���Ӑ�׮�����e$��q@)N/*��(��3��l4���D�J�DE�
��8Y�TÅ؜��W�c:���,��bCd�ۣA�	le�(9���t�����Z)�OnG�O����+�)�j킳_[�����#��zwI�cT"m�v=rG8�=�8��(���~Z ����V���H0���%y�ם�M���F��]��h]��.b�d2yl�){�h�
gOT_�a�h@Q!|�p|��tG���[U�l6��mU�Y�ڶ�_����~������u��\�;�ղz؈�x:��|N���}E��_��</����ն���MM�W��}柙��9~cU҅���e5�|����V)]P�].��ݖ]ڼ�q���\:G&��"+�o9*}*\.w:��LPM1,�
�W��c���*�u��ܕV*:���������G͵�X���!�ae�N�c�r�,J�5��N\\.�m,)D��@�E>L[�w]�27�	T�ʉo*"�)�_gma��7<��o�]�j��E�|lwYi��l-=�12r�ϸT���r�U���]YXB�̘P��E܇&�۸��;�#g�'L���P��Q�&�3�_9�}]�|�:B�FK��$���59|�X��wc_e]�+�N\���\�uEw�"�r�Qsz͞wL��ڛm0�k/v<��Ԣ_c��wÜg~��,|��2>=v.����:J��g];�~3}���EoG�3w~mt��GF]�l]S����阤���;M�Σ�l\���4M�l�Sw���d��ģ��v�k��� ���2�ov�ŵ�4o�b�ueo|���5�'�xp�v�,��9�Ö,�t�!�5b���P}Ovx���b��0@�r<+��<���p��/���j��1y*�>/��k܇3�8n3}�qi��WZ���b�~��}ǫ�����`���m:�t_�2��߾?R�|q]B��A��Ѭ0�8����Z���z�Tt�|����(���1�xE�Y���6��vRWg��=2��E�z���ڇ�P����[���ԥmX�w|O��u����Ȯ|�O�S�+��҈��U`�l�*k8���c���h%�@n�(����g����q���]���c��1[�0�Rf'�B�8B�.Fx��-�&���]�A;E�~�  L�i{�����׋4��8��/*�v����,�mb.7my�ۭ�����I`�/��fTy@���t�΢a�/Du�sj�*U���Q�7��J�0��=f��g1�
M�ӨI�r�I(E"w�Γ^p�Xo�y.PTv��J�R5��:�)��� ], {��3�^� �0���FT�;�Sxr�v))M���aX�s��E�\�mNp�Z�y@=�`�\�>�.<mb_vE[x����
պ�6�\�E��;��`5H���O�dtlnp�Qc$2��U��[7
]�5+ێa�]2��|u�9�F"�Sb�G��;�����v��^{���/����g��;�d��c,SllШ&�=À�1ݘP��l ��0ipG@H�Ћ(.�����<;w��汢'�h������B�%�K�U]m���>���N�FB��X�k-Һ����,�S��ũ5Ӡ�Qr�2_��Ճ1`9S`M��I�!�WU_&�c@�V��#.0���Z:�X>K8Gצ�o^u)RQ��Ļ҂˂*���p��6�bq)��>�qx˦�����f����v��*�׼�3V��C��
��v���hM�8�����xE7�z�w�'U�	�׫�P��'!�����7ِ�w!ƾ2QD�ݻ$d��Li.okϵ��Pxiٺ�gF�ꄌe�e����jQ5�f���f�,�a�N	ƃ�ξcR��׋�r�kz�N���``r���dxH��st���� ,ӵz�i���;�"��K�i{�p��L;aM<ј�r�Z����|���O��p�:�\<�zs��܌Ƥ�(&�N��e?[��$�6b0�Z���3���̾��=���JH8�v�������T��z:�r=oг(������.���� xL'��_+�	;�b�?�)�T;�!������ԏ�OߝNy��
xU#���zl�"��(��lΉA��2	3��@6/�.�&�خ����{�2�}�k^��y���A���`��F��U?��m��ۊ
��%gS�z���Af;?�"V��P�6˖	�	3W���Y���N��/?5�H·��j9r6k��D�2!��H�!<�.|yx垼�Ҫ��ߢʫ�t���q���Al��\�c�Kr��Nz�f
��%j-r�U��+ �=FӍ��"�qDp)F����UqV�' ��~.}�v�,Qe,������RT�(�[9r`;93v���K �AU��-2��H�$WD,A��S{Ú�=��R[B�f�S�f�j
�g��}�ڻQٌ�&5��TƤ�n�Qg��3b
"��E3�s`_��?Wi�z�nO�L����?��y�z�^�����s���z6�������k��1�׽z�%�6|ާ���$�Ѩk��*\���_I�[nmU�
��4̊��
1���UP`�
Ȱb1E��X�&n��D�S+ɔj� � <�� �����c��=��{�>IE�oGR�C�����}6R���|�k��o�������l�g������3�~4��Y�깐�"� ά˛~>��������e����w~6e���e�R����h�cdߍ23'?��ù��j���g����O=���-L�SB �2��
���!��n�bˇ}�] �5���<��;�`����m"��#S>I��X�3 ��ˈ���gG���4��lչ:ҶtS��fl���zR��(�+B��qv��Q�i�����X��/���L���d\y�(���(#s1_�;����w��Si��d�(�ݗk[�K��-�b�|3��4�ޑ��*Iڐ�r	l���
�J|�Ff��E�^��bT�D�b;󝅮S~CM����2=&�F�+��X4�貉�֦yLk���)q�P�ױ�%�j��V��r�1�trS�����$Y5}t���a���v�#��]L:����,z"�u�Sr'a�;w�u!��SQ=+
����씉(�hx���y�͘�	o����_5���u���JL��9����������\爦�0�l��8��(ˀNk�j�-9�àj�N���%a8�@��}�, .��yޑl+<����f�\x�|(� �	b�����b�'YB�4A~�p�u�uj��Tũ۫�+�N�2&�A�%�E�~s�����N'�����!�w�>>,�ޒ��$d �`�)� +�b	׶�� ��m�J=�ʂ@v�O���4ԹǶ��ZH(���T�B��|I���/�̏E�SA�K�6صZ��,��%����a�+�ߩ2���.��]3���/���4�Z����l�Jr����ڒ8	L̨"
c��a����#B��Y[ij�Q��!>�ޑ�s����˟P�/�@�B�>�eU���*C�\�)��l����[��F��Q��9|�>���K�3^n&� N)�E'O�$a��|x�YR�kan1D�>@�2�����FR�RkK�Xo�؜��%�20�V�#�0<O��6.gj�[ߌd+�{�<3�ŻIy97�f�A��A�s��pa/,�� >�u�[D�kWOt�R[x�B9��zK�V�`� l��Q�8�.� �h/*�n�椝%)�Xʻ�IDc\IÍ��rq�kp��B"E�H2py�_��<e9))U:�M%�hv�kL`��K�Rȡ�--�H@�1�u)_p�V!9�IW������T��d`���0�{l����BT������@��4|�o7Ț-��{r��Mst&s��' �:9Y��C'H��F[�"g�``i�[�a4K��A&�}��k�g��T���lh8��M�O1��@�Bu'u���V8I�Z��pjXiy6w�Lͪ���P%�Y��!b��"��F-�a:�e��;G���Ҷ�y�-OR��Yy�LW�m@�;���Cj@�ke6 '�R��,��B`01ܗ� �4���o��#rufR�(>� A!?�O�삤�U�C�B�ّ��p��sy�o��o��˾��7�zߨ�}ޫ�ڻ/�sS���z�g����n���@�6,����ku�)Ug�)��Ϧ�q-3���*:Ob|��ɨ�;J��o
��8ך����$�1ӭ^D�n�=�ӱ��&v��gmN��3u40*����g�vTv8�{3|��n-t�xM�)CE+�����/bJ���qu2�5��C�A��3��ԥo^-ѕ�t#�l�T�2I\�ݜS1�l�\Oj�/j��ۗ���Jj{&QLB;�2(��c�5s��#���R�`��&��ױ�B{T\���<�'+����b�����Ku*��iױmM�T1TV�����lL]�P�Sg_A�����zی��O�9��27$j��wU��Eͼ#&(�La����\&�jу�I�*��`�GUa�:-dX��"�i�G&r�eVL�2������X9����ց�n��jz�-]��讝We}fkni��ܞ�N�v�dt��u�q^�6���;I�1�"����s㧵��cr��vcml�c"�韙'e�iՆ��oHQ�`���V��)�g5�NJ]}=ݥ+�Ӷ�؊lP��+6Z�w�{�h�.wnqjk�R�w�
��=�<r�7��3dH��h��7{C[�")_q�h��%�.���>�z��ȗ�P7Rw�5o��g:r'��?�p/t���-����NkDqUE���ȥ�;R�[��u3ׂ��*H��0��ɀT��ʍ���m�}*r���v��3�E	�h����aEѻ��O�,ůWZ��*w���ϪьP���:w�W(��N8�[���瘜�k' �%�d�H�=�!�uؼ���#Oe��)|��GN�OV�)���XF��u3��3.M�t�/P��q�0�\-�c�;lՆl%Q�"F��v��o�2c�;�2R��F��˭�ѱ��!9�LY��G_R�˦��.�p�Q��5y��J�fnhe:띘�ULa'�r�[��׊nF�^�T�����M�]����l��rj6"\L���{sN8�����YN�H܎���ML#�b���DS�>f\�b���=UʇS�4)ͻ=y����frp-o3l��Ӻ�]|gn�T��d|f�M��/E��{�6~�$��j����ܬ0D'w��_�6�]FqCq�@�є�FՅQ|����i
;�	�w=��fE'ωym!chS���1]�,6
����{3��6Ɏ+7c�/���.�c�.p˭��y;ʻ�m��J�ܶ����yc��Юr�s���g_IjJjJ�xc�w#vr6�L�]ZMV�.eN�ȣ�uAGu��K+����,Y'j#k��fU��E+-.�CI�r&�$��;
����H,q}��<".H�����U�D�Y�&�x�(��ط3n�c*��#�\W9Ro(ʺ�3�	��D�w
w*�����hefۋS��VwҾ���:�s۵]{����[.��}3��=�I����v�]4DX蒢}&n����-�2u�a7� ��uY�X���]G���u{�Ce�e͛�i-�n�`�oU�Q����?5OϒP�����rev��78�8��yg,�Aƺ9;��Ӭu�V�(Rr5��B��ɩĪbc�$�o��������1o%�t�u)�T��Vj۶�Ep�ٵ��6�|�vRu�y��Y�|� ���m�g��W�3���y�{���I��9����y^����	5����rY0MetC��U�f�e��F>�[V��Ί�wR�	3��֭�B��M�Ⱦ�NM�����ź����N���'U��[��E�r����;;v��W�W{V\�Mn��*���ٹ��Pc*2.'(�����ڤ���u�c�mk��J����Nt�2�g^�ʳ���F;l��1�Q}V�,�g"�v_�&c'3L�R�r��6��;���wN�L*��6b�RԷvņ�)B��pCY�tV.L�ʅq<������d#��n#\-�ɾo�����wz�Q;+c5[�ʹ�↥�`I�vz��\�lQz��A�����SS�4kA���"E30�%�VeN�� H�(<4����û�[~F�)�iH��s��-�PΗ���_A������������7�8a�mmXj-�t�0e�3z`L�yA.�릡-���^��Q�9ى�Q�����y�����f�r�%���.��G�m���fnr�]T��MÓ�z!���7
��)�U�;�|ܵLe�)�\��B"6�Y7o���jU9��I}K�d��n2��&DC�����4D��]�D�TQ�tH��P8�Rqq�]@��v�f[2#&1과���;��8�ɚg/b9�{E�s�����\ٛx�w8:ȗ2l�F�Uӈ��=�&+��
2L��u,x�{U]��#GY��E��Tix�Q�|�ou���'��P���ou3�M�D��Ǆ&hW"�R��c�ܔ�K��<�B������T�U�H89f`���7�:��ؤ�
�>�l΋�!eڒ ���YBr8d��S��=+�����X��N0h�u;�*Zu�V���5��0p��\�o'"&y�%���>du�^�����|꜇r�8b�1�K�[�����l�P���"�<����n�k��G!s��H�x��uE]���"*����+���݋m��e�5Ze�2����̉��ǵ��y��|65п��A�댣JL-����j1�L�7ƻoV±�:H�&gA��<�'#s�h��1Oo6�2��ܺ�o�	7�S�f޶�&��9q7=B��f�����{�,5��L���U����\օ��q�X��Ô@ݨy�f=��~�99�yY��W�51�3�����!7B%\�@�{=pN��)!�;�����ȅ�M�1<ȸ��:�+�-������+y�C-�QtU'�'�6��ۨܚ��tj���4����UU�js*U��D���ʹ�����Y�����7��R�ڻ��:��s	5���~7|on��<�U�j�q9
R�F���w>e��f,IS���E�֥�w<�F8H��Ww4�%��r}J�a���S�Dc&�ݾ���a�8�vuɪ��ɝ2Z��D��Rv���˘��u�uN3.3]u����1,ۗU5*k�ͧt禺�e�V� ����u5���2ud�sU;�W�H�����: e����f�梴Z�rv*"����+n�:o/�.`�5��)��X�"DglI��F�����ȷ:-���"�v%�ˎE�K��Д�u�xYV��9��if,l7ܡdIsH���(�{p�W=��T�[+��z
zaPմoj�.����/N
/E<�f�'J��t0�"M#:n��f7}�:�e�k�9r���5RH̪}Oz��j�7J�ީ��7Jv��2�)�ɜ\�����P���l+��f|��Y������aGzD������F{0����g;��k�{g"\�zN�oM�g-Ȉ*H7�1T'o>o��8|��U�������v:�/j"g��:���ٝf����X���e�̺�7܎V�B�='�<ڻ�33}ڬO�M��֬s��bRv��*Ę�r�q�O"d�c�Q�L��K��80V�U�f�f�A]��1��4J��͹��uiV��u\�2�\/}x���È�7)�'1�L���2@��}/x؉P�� jF�L.��7��AA%(K��|�(�K�˵T�C�69�F��q�6�{��q�Z�3�;���B�:�SP��W"E^�Ȓ]���8����h�n�qr�����\�z2w�m��Cu]^n�8p*�_b����gN䤰�^�t����c]�rݧ"S�=V��o31�m'��%wu���7T�A���;�|6�f�:���[sk&Ӭ�Vnƨ��Y䗙�-H��8c��	�4�%NT��՜}4��nhq�ĜSѝ=.�^S���ktZ�wZK����3�ć`���	���YZ�r˪u,�G�\���F�8����VN�ou����72{ \��9�Ԫ�{����7rA�V2���7[��^�	&�y:<^�܍�1*�	���ͱ9�j[�Q�d1���97FV����Aq1����DK������VU��X3f���l&,��|�͊ݦ�l���)��gL�힜5�y52ui�x�{T�<����`Q�����V�&RC2�n-�"g�p�N�"�f�X�����&"�D�U�]QW��ڂ�aG8�G��v[��j�w'_w4���G@�'$tQ$΍;�H���.ɸxc
�*&�p����Uz�}Z�m���GgV�;;әld�sF�2V�ފ����%H�۽)i��9�(|�PL|t��ع�Cpɷ�[��{�y-�Gz1�d�]k.I���{7��BY.���3�>q]4*��Y5Ѷn_x����սw#w5�p��#�P�X��4�j����Φ4uΓkOoj>]=F��c���OB�6�q����L	����J=������i�݌��p2+-�5MP���q���<�����Xo1Da��t�TJ-9}c6��0b��@���[ٖr5dJ����u�W��3F��������l��L`Sp��f��GwVB�+A�&DJ�{��;+�&��KšS�6z����Z7mV+�+�y�R�E�F��H���k�׫��YH\�+R��&��[�&���9�:s&��MD�Z����{q�3�����a��2��Ы�[4 -�Cܝq�\�[8-lޓ�:蚸��#rz�*Y�S���Cq�����+g/͋� ��ɒz�0�t�F�Zڮq�<�2�,gJ
{��fB;q����仺n3��wJH����-[w�á������غ{���`""�l�m����xE�-{{��I�� ���u�����-�5�h]����S�3�U��@=���p�)�>e�w�*�=3{nFJN����޾�$��7E�d`�Z�6��Vq$��],��1��A13�^>O'�e�0;�b'lG��بν��͘�=���jӱѷv=y7%S���U��T����^t詭z�iS�/1��M�;e'���ؕ:���YJ(A��m���ĳl���z,X���x�s]1]�3���%t�k#*��z�\�[�}�oFO	�!��*����f����X�g�j�ڻ��9��ꩉ��N���yu� �����Ř�h���d�C���GzL���ne�A�%�S�!�鷵�{s�䫫ۼ��9}�<�,�͈l��RF�u�KGK�F���+r��Zx�p�.���t2��'-T�ض"�f⃥Y=X�l��r�^�E]i�5�M�X���Z�t0N8���d�%���za��!��;��ݙ�s��;��_gM2�Nv�R[�Dk��"�#��P�1�6��.���n�9�O��Uw�;aC�yfc&wxnᾂ��MwJӗ)�/N�K��v�T�ԾR�l�ˤEWSΨ������Sި���m`�W����3�T�Y]Q�v�c)v9w5eݵ	�i�2��b��YS�8Dl���?-u�ï.F��[�3�鏗S;e��w�ԧ��O�v��ɮ���5���+/G#fb��t3_D�TJ��jSW<�jh���;ö>R B��u�QB�C����*�Ţ�t������{n���;��*���bcHʍg����uB�9)�ˎ �E��*'G�^�!:.&sq5�M��Q�Tl�WTֲ����Pr�I�w����,�Uo�1׏^���p���ٙ�����q�D�nET�P؊�u]���l��Q�i��v�F�]5�������E���|��/��,پ����u��o0�Յ�|�VVsf�F��������#�龼�"l�Yw{5�tvY�I,�U�6ʛ��g����K�]�h�p�st�U�:��,�T�#ض�w�\\��Z�kFF	����,��u@�q�@�#M_u���Z�98F�Υ�Z�2\�=�W$��TT*.��s���8�'��t�U��g.������=m�m�7�эnh��(O.(Β72����;�;��y������L���o���gRY��f��?6_3�%���/�b�'��ɩU�.�υh�qO6���kf'����8۪�z9LeLqX81ö��|oa�Q�"��d����6S����-c�싳VcV�R���f�mt�;�cǻ�#9U���ntc��|�T�j��rQ΄�g(�fL)r�B�LH+.��a��&pL�
or�<�顲2��n�`��34vR�Q#�3L8��G�
U�6� gWVrx-�v���ѵB�a=����#�_Y��F�D)EU�|�Y���LU�/�ksbTǺOJ"��>.���tRގڈ��d�l���7�,�qj�o]2:��\��b �s" DŹ2�o/M��ډnb����:��T�P�c2b�\���ŕ���")[] ����[��VG�I�K��kVT94��Ї���T��tj�ʝ먁;�'n���#D�eu�௎l��ឹ��'v�w^�mƚ�#z�Z��X���բ'smQ���.��������mj��1G�$��1ї�-'�D�@�$2��9�1j��p黧`�v
NE�'s�f��zM�<ګ�4��.���3)ED�����1����������$N�S��,|lN����ک�����ғWԲ9��M\U�b���nb*8u�g��B��q���`�w�{+��/nH�yOU�P�®f�Rܓ����Nf��j+�U]��[�s�gN��0�=��Hw�5q�Z�W��*r���l��[�n���5��ݔ�K��y����귍mp�y��;7��U;�eD÷NY��׆w���r���蝭u�j�V�l���7����uQo�b39��]!@1��*�=�l�ڷ�*ǜ(N����ݷ0�Z�T#e"�&{��~T�����P�wF��X#Q�ZTX�kjZ��M��l�V�`�Z�QVؠV�j��\��,ɵsŵ[Vh,�!T�!l��,��%I@�,�J���J*�� �,d�#�K*�"�*QbҴ���eU�ml�����[&ckFՇ4�f�66�F�h�V�)m*��EdJ�E+,E�������V��E�������eJ�ƥEU����
�նѴ�"�-e[clZ%b�j�`��U�U5b2�(T-(�P�EB,*)E��ld��*ūJ,m+-�+Q�,��ִj0e�-�K"�kFт�Q�[Dm-K�*%F�k-+Rʕ("V���U�YR�UYbԭQ��Ym�K*(�ԥ�`��+J�H�EEP����T�e��"[kU��*T��j*��EQb��UF�6���TV[V�"ȭh�U�--�QT,Q��j���V(���R"�QQb�4�FVTh���Qh�Tei,��U�j5��I	I)J�l�- ��%Sv��]�]��-��[�~�ތO���� w�.`�ߙ${�W�=߱����}��]�8CS��p©�((r<�A�~ ���p2����|_�=�?��Q���&`#��$�7���c��#�گ��S�׽���.l7���r�S�|"�Q^��ë��q�Zc�_c��~����pg�EF"��1�e�祭�u��<�������F#4yl��#��qOZwK�"�k��Zf��	�Y8MʟlGo$~�`F�^f�,�O��Y�.K�9�s|�YW��X���^�u��"O���+�goz[��w!�.���mJ�W�����ϳH������^�����v��<b�޼o޵,�3=3@�*�5��Ь�c�Ac�gX�zwV"�F��)�ÜL�2Tz�y�4�1�[\,��W�{��"����t��F�����@j�"KN�wf�[�9�f�l��)�]|uZ<,�a��E�X �I;q`�.�ѫM���Vx��p�Or�q�d�1���$4ܬ�&!9ȃ���A\��:e�s�C:{�i�yrMQ���nf#�U�I8+��v�,}������N�[`����=
I2��V�8�t��|����5G���L��c���t�>q�uC��,]p�� �����{3��=zHS� �7��]2��ڊ�cq�>��}��[j&,J������ �yml��é�T�c�{_�`���	�!W̨i=ˉ�؊$�[�6-k�mn�Q:#����1�*������N���DoXʋ�s@V�$�����'F���%;:�s)&a�'�`�-	n0��Wڰ)�G�~�F!O��v����gp@ؖ���\������W���P/�M-��i���A���X`���$-TZ��O��R�T�����%�:z`\��dQth�K�:k�~ULːL��z����PLI��6Gy�W�.\(�BgS��K5h�J�r�8$[��1��ͯZ\����9�L�/��s6*���Ѡ}r����뾗:��͙��edq�tZ=(z�<�����h)b1�q���Ϙ���!N��܇�ڡ��;Ly�<9�d���Uܔ{�\��ݪE��[R�)9R +:�[�A����q5���$��j�V����  ��yw����{�#�0+#�!I#�����C��+��?������1;�o�O��
rD
��A�Y|z��n�&�`�Y[�K�QG����߃�RPx��4ObҬ�s�SJ� fs��Ƹ�M�kcKd"���aAD�C�-�~Ì���q�PhS��v���j0�҉G"�����A ��J����s�t)(`8��c:23��r�gJQ-k����Kd�2��(R�c
N9<�DDξj�$2��q=�S28BRbP��k��u�Ft<��*MR�RkcR��"QHŦ1N��Y�����e��$ �D���r�d�~�]�g�w{߇����K�ؾ�������:k���:L�Ӳv�����5�Q�qtA
�Z��/2T��V��^��S�����zн��{��r_o�=�����"���Z7�(��KҠ_�_̀�A�}�}��j5	�i���G�< ��E:j�������^��=���!O�PB�w�{�|��Q_�X:��-hϟ���!{�֖�6���0w��ΖԢ�q	�8�v�x  ��8X�Ӈ���ynlu�6{�y�`~�����%c��1�2n�GX�Ni[3>m1�!p�Q�2A�F{�<������������뼞�w"Rx֌h�+�'��Y�ni��2ѿ�C���g�	�)\F�V�<��+ofk�i��1ﮑͷ� NcZ�a��#�h��A�5� �GO��2��{=�K
���[Y����p�Y^��v�0|yMPKn��!-��W�לJ�_2CY| �<��z)��N�v�^.��a�F�9Y=Ӟ��@tu׿H�WyԖ��n&B�����q�H|�xV�y���j�R��ӣ�vh�_�5g�<-���kO3���v84Kq,s",��˗����N��Hq.H�*�T����r��n�E��tv��	4qKʓVf�w�I�l��6�i�ՠ	T�:�����q�0Z�2N��v	��cC5D+���x�>MO6�S��n��.r�`f�Ɋo89;s#����Z3W��!���DM�Aݘ2#1v�;�|�ݱ�"��E|0f'�z*��E��EU��ϟ�;h�k���a�,���[�+�mu�V}o^K�_+��RD�'̪�����!��ؽ���6��
:���l�:h�XD�G��X)��3�Ǥ[�,VQj�޾{�P���Ց�GHC�%�y��Z�)D��Z��ǝ�"��C:H�]�d�\�Hrev��d+��ˑq�JݟT�hP�2�#���;>s�
��0���*�U���+p�y�5{�.��$|.�Pp"��sT]kRʣH4��8o�)e��S����!%V��H�~��ʭ�A˟Ö�<\�S�G�EV�=�!{�]�]��5��_Sq|v'��Mmp�U�G���Σ|�6������(m��&Ew9�i֢�2����V7���~ܩo�S�*͠���+�и��tKe�讼��u�7�G7�N��Q ��/zm!5��}�,�07As����c���9IFn�n)ȯʾ�l:<�5���.��m����vo�4v���������VVYeu�PPz�T8�Ҳ�Ì�e폳��C?_t�7����)�\,�������	\�YSYM�8اHL,iੴ��1�9N*�f��� � �@��ԣ|�lB%k��"�J2)e+̃�1�t�9�1$B� ��T�	�A�:¥\�zK#�؛��i2���O�jbIte�`[X5H��U�:�x@X���|��-˗11q1���.���d�X�o�DaB"�R�l����Q1�������\��Y�;֣��}����9����w}[��:/��}�������v?���|�{��qs����>�;E�(Ϭܫ��8kH�	!	F��]�W�hu�w_����l�*����H�A��Q�o�>�r�~�t�T�2����C�f��/z��+)1��2��P�H=�*]D0Q+�Ye�bJ�2�G89zZ*b�e����(��R�k�Ka��)J6K
Y�"u ��*Qjb��R���s �&��j슌-I]a+�0IC*Q�y3bL�(��D�+Sf�'����<<<C#��/���څ�]��A;mK�����_'���?w��5m�������ղ�?��w���9l
���I��Ogo����몮���A��zUH�꙲��3#[i�lͳi�.���bd�bj�L��Q�E�RB����4���d+����I\����/^�n�����|�_�����_}�!�	2TqF#Ƨ۔�}^��i�? ���_U�5_M�+�ܛ�;AQ>�}s�A3~�ٿ>T���2��F7�e(��;�ڸ�ϩ�����e}b��}Q]��oOt��LuS~��1�V��<6�h�~s����qz��}��������������}O��'���S����~���O���|< |�����J�SP�}���a�#�/����N@��-�����pk�O���i�n�Y~j"�z8��**!*ڃN�.��"�J�ov�*�h�[:��)����W�w���I`�����	4I6)�����ٟ3��z�����nOs�;����^ow�6�G����;/׼c�7+����8��������Ѫiz-�)a6;�JB�*fˎ�g	O곶�74��׆�r����|������C��n_�({�g�,�.aV1[���0ͤ,,�Yz�����m����:;�\��<q����;'q��O}��+���q�?PU[cȏ~�!��|xo�����z������{��~}`<Op���P-�<�3l��)�"{g�9�>^���m�=6@��������X��O$;�'hO��N��z��F».޴m���K���B�+�s�����������|�=���:p~��N{�����a��`{ho���;:���5 U��a����LN�
�K�0�Ĭ
��l��,p��Q���Z��)@�v��:�c^-q�,8��00ppm�n\d�?����+"��D�����Hd���M��S���)'���4'�2L!�}�i'�Ɔ��7�]І��ē�^>쁩��O�$�����ǹ��$��	g���'��zx�O����z(�����'�՛�x�E`�0�֗JR�H��20�$�߿�$4�$��?s�~ϒk���()-,`ɡ�1v���*�F�ֱٸg��r`���Em(2|��*��V|�U����|'��{�1&3E�,���1DW�j��{ek��+4��QDI���-��m?Fj)�j�0���OPɌU����\ɷ���R�-�m~����r��b��d��jD��Ka��4TFs�K����9��b�N�>��NV)�/�n��QW�����*~o�7-��J��-��3o��{���)DAJ�T�b����dTtA����V�62w�����ު�9�C��EQ���UX���\'qU�����矖_?
U<Sy,��y�����⋠���b`�ڕ�����Y����D#�/"Q$��B_ -݂/�A��?�Vq�j�)�=��Jʪ>�N����G���B�Ɗ��h�Cv�v�QW��ܪ�:���̻�v���1n��w�X�����#������q�b�L_�T(���+�?}l�A�I;~�ŏ�Wh�Q�)GEr��-V߾���N|�
�}FG�?��>���a��|[_��{��^���=C؞�Qm��{ʶ��D��.;��j�.�3ǋ=�����i�=��ֿ�H"��Ϫ��~%a�v��������涕�,>>����%���N�;ER�8��NN>D����rX���v*��� ���}{`�p��
����-jT�|l������7��w�ώ����"�HI%LHa�J��~�a��&1����R4�$<�>���;�C"+�LD�RI I'6���y�:>�q�F������y>Y�
!�����g-�l�T_{������{���u�7��¶�h_/߼w���}�{��5jk���a���,�ǟ㼢Ҡ�|������->��2h�[���~�Au`ڏ�͌�?G����Ź	a@�
m���6�?���z�bۿ����iWة�Y_��������{�F�4�y?A(���d��ñ�[@��*2�O�����{��������S�88mM?_c﯇ɲ�Dx��߷��	��y���Q�	!��������-�5�?%�?�=;�e���6hUE�:<yg�}���{��W��e�� n�Q ב;���,a����K�o֛�R�����ض��9���!q�!G�� |J�1�IY͗K+h��Ǒ��0Q�Ɵ�z�,J=�߼'׾H����{Ǿ6Z��/oD�*��\�FN~��}�ϡ�*�� ���� W���g�{Q �K_�rM��P(�o�3��� JA�Z����>t;T�NO����)��"|b[~�M;Jҿy�||���D/zݳ~H H%2"P@���-�aj�Y��w����Md���J))f���Wx��
p~���Ԫ4��>��겠�{�?��Ǽ�ZSϏ����(|Z�T7t1��~/׏C<X���2��W��
�A��?���8!��l�� �M1M��K�k
M��|>�jƾ�鯏C"��O�����O�[ꅉ?O���^{�9���@vS|�P�
��Ay#�nػ R[����-���8�1��|>̃�HB	�i+w�x�x����	 }b׋Kv1��K� 1��>|���)K��0��-W�=���OUs�����{�g�>xO�����j����$�Ea�� �����BǮ%R��̓1e�~�&ÏR�����?zHg�{e�*�d]� Y���8�ݱ�p~�$`��0��4w?��U��zA��y���@[���C`Q���~��6"�)_}���ia�y��9#5M����#;��y��%/��5��;�8x��Z���>�UH?~ 0��O�t>��	�2�~x0|�p~����l�/��Tm����H ��D����7< %;�s�*w����9�ޝ��a���a)Ӓwa�9��?g���>o�~�����~��Nm`����C���#>?���'����
H�J	ac��b�c�-����^�A?����������8��m��$�$�Kl�-Omp.�\�mK[,�1�`�x���a0\�3CC��a �C�Gn����c��J�;���x?���??���|���G]{���x�R����zH���z[����{�ā��� �_n�u�߉�ޡM��!��^8�OzK�t��Bˢ��W����O��ǡ��O��EL��=�$L#���`z���ط����>��q����CS�`����	"��W�f�@�,[�P>ʣ@U{OdǂX�߇
`o|�{�>7g�x`�Mg�?=���gl�q>{AI�����fB&8/�x��oC��L�x���� 8�\�ā7�[�I��o,z�g�X�&�z�O��<='�};�6~ ��뻱�����׭������nV65�[��v`�ِ�`�;�� n��߳�π!�_/O�d?)( {�>�����.~�v�� (ܘ>�=�O'�<:��|���O��~����a����@���O��dne˗�"�#a�h�Z��cs��b�}��S��/�00'1~�� 0�)&L	���4�����({ۡ������}:_FCX�`|u �O��`k&L>����N�?]��������|���.����?	��d&a0Ʉ�����O���������'��f�P���=�4ӺN!��L!��?���{�w/K��)��t�]t�ҝyXCL���W�N��2KI�~��Y��G���x�L��'}f"I���B��L��h�%;?�Т,'���uDTs�*��6m	~��i��G�x��~���>��Qnf
�u*�����+>�f͋�4��NDb��a�Õ��,7M6m�i��EVZ��,;��QVQE@��$��D�}h��a��'�r|�X*>����֪	������*�qO���-^����~Z����*)�*ݺ�m���>���*��/��2��[��3�EDU���
��<g��N>~8��D�2�Ҷ.L=���S�m8�s�O� ���*�l�Du�AUuG�:説Uߝ���F�R��������_�����^F*;�L����X/��08V`�����ȣ��K)��Uɲ����󦚿Vi�aZ�D�᭑��)���<'�m[g�Ӷ*0]�=��+0Ū֕O�=�ڶ����h��qꭩ��e�����'x��5C�+-�N�O�e�O[��j5���vyR�������mjW���0Q�<�J-�W"i��=���|��zn� ����wϻ�[Q秼���T�̘UQS
fҎ��^�b�3�``E"~��+��&~�����}�>W���*�����Af�G�w�hÓ�B�>�Ͽ'��Ջ�_�Ǎ�%F(��,�����QU0����Y��+Fo3���ʍ���wK�m*ң=qا��ߟ)_�<{U����j��������pX�v���׽���JS���+_y�o����G�����V��{}Yx,�u��D�R���AD`�p��p��5tܭ���/���(<{�>�>Iw�M��ez�}=��	 	wm����o�F��"BH	'�[M�E��q�>Z��w���Dy�i�|�`�
 ��h��$
>N�����	(���K4Y�b$ �K��--Yih���b�K��#�������I"	E1��o��ѱ� �[�$�%��Q�|U}��lU�������#b�"<���b��"�$��+��C"o��q
�I���R$��L]�i�H?|�~h�4���$�s�b�ٴW�>��d��A �}�~�}��;�V�����;�(��ٺV��_��q��֩������ac�W˻!7e�4&��W���n͉�|�O"���P�G�����ϖU^�^�����+K|{��/��~(������O"��Y=?_�O����O���v�������v$���D"(���n�hR}��s�%/�+�&�N~����-�>��w���ק�)W�����i�>���Ų���ӄ�S������/+�����P�,~Qӌ�:���k'�{z�V�T{�}����#��{ͥ=)�E[e}S�������g���d���J& xX�3�V/؄@��6؄H@��6�A'�:�=�0�}4f������NY�z)荟_>��@�#�w�>�{���ڥ��S�C��_Ǭ>
���è��m�����x�H���}'҂	䆲w3	�M��2Ae 7_���A%?:۱�Y	F�
������E���9�g��~~�w�	�a�}�v���>�ͪ+G����W��i~����z���b��i�-=���RǾ{��c��@~;���~����K�}>��y�3*Q�̻����e��a��$z#�W���x�C�ï���ϩ�- �g���zP+h��l���G�{���wbɼ��>���`U,�Ϯ0�Kb��ނ�d�D�t���W�����#yb�2|׉^(�>|��~�>�F�Q��ow��x�����]z��b� ��n�d$
"A���f�<����
g����(
$~Ü{�'����ȤyC���C/��~?��$�x�1S���:�	o�I�(247�Mx$O��X�x_���l^Ե�Ǆ��ߍ���/��E��B�ף2������?DY�����������PN3M��KZ}}|�|���w�@C��_>'�԰��t�6S��ɪ=M�͂�n�F�OJ}�;�F}d�$���?���y��8�Y�pv�2��~�&��zn��������g}���OS�p�@y��b��5"�q�����Ph��}O�<NKj��������pٗ����c�Mx��,ߘ�'���������o2/����tx�)x|�Q��"�>;c������	�$q{쿷=�h�j���ݗ�2 �X�{�e���"�����s���<���!޲2�S���� ~���~���I�w凳��l��>zrC�~��.Ņt'� ����~!����z������|_x��y��!N42M{�u��~�6~Ot�qR�~=4�=bi���=���ʧ�zo΅g��z0^����y�|#�Hq�h��� `����zC��x����������������f�8&�;��z�y��}x�����%��e��HRп%X�t�D�����0L�0�+-(L��V�ʪ��Z��F�|^O��ֳr��n5�t��%;"�����[|����;�JZ���~'��{��O��R|���2Z�+Q��i14�ZMS�~h�t+����s��;��\��d�_3X�� *E��|#L��Y�m
3W����֡�5����O����>8*�}����Q0X
c������V�"_H�A�*@<n�zC��aqD.1\���f��q@���XM�+ST�jM�l�^�Z%B��}�����#yJ"�����Q㷢Ĵ@���;�X6�
B�b��@7�V�B O_�4�U�;�b��8�Zh�dqS��M���8��.cd�!h�sh�I-& 2P��@b8,�Y�M�ʏ�i�6;m3r�) V �)+r�Lap��[J���Z�>.�x�E,T� �r�d�M+)�Q� $�\�Ħ+U�WZ�|���-!3:^ϭk`��w�\߁�Uj�s�gGo��)��	��'�:�KU�0@K�g��1��|�a�@1;˰~�i����q@�@E6'S2�ɧ�lR�yO?��?f�q��?��!78���=��q���N/����B �0��{��d��.�;�{{��a�˽�u������O��4?j�-E0b�X����Gf�^ʂ��p�m}��;Q�!��|p��[���O�#��y:n[�;��<�C��rV;ߩ��壟�.7=J��:ss����Q5:^�m�f%��:�ڊ��"m?+���/FC��x����/�]�ch?�� T:���3�ܩ/���M�/V����j�C����D��[v�s�+z �H�ﯾ*T������a�n6�wZK�������|�P*+���_3���Yr�8�W�$���
����5
�"�Z�g�k�w
7W�~�<�.o��Y}�O�F������6oݒ��~WE�[��I ��o����0;���o/K���קg��	^��.$���������}�6�Y�R�cADF@��F*�`-e���J"*�-J��*�dV�$�����"���EV[E�*��UH��h��[6��Vk4mL�,UH1��b�� ,X��$���S��k_�r����;M�`��X��\�J$bKi���9����Э[Qk����� ��b�9���R����� �BB�>|"��>�>\_��e2�mKs"�iF�wFj�n)��Իݨ���V6�vLSjf-�A�&�M�� ���{6lٳT���2d뮶Ǆ��0�V(cP�e�����µ�33 �d�`�2A�̔U���E���,em�m��
Ŵ�"�=$�!l7KiUjV,X)F���kUmPX�R���ڠ��*��j-�Z�����32���T-��E
�-AQX
"V��(B��Z�!hڲ��@����%j��ZTERҲKB�,+R
VV�����j��[T�kF(�ұB)J�I)
JB��q���LJn�M�Pp�|�?��⿮S�re��������MT��7���_�֋ݹ��,��+[��(�Qq��bV���n"Z�Uʔ��-����s��8�2�n1k��L
k.��b6�AJ��Tƈ���Zc�����s-��̣ ?�'�1����]H%Ab�����>! *�`��z�V+a
@�M&R²��b�"��H=�-j�)[KT���Ғ�1-��J� $���,7z��2�l�T��4h�K[J�-*[RƔ�V��?�O��t�����i������_����0?y�>�ّ̹����u*�m�g��WF]�I����S[R��O��0��O���4�s�(��ef#U2�8����������0)j��21QAH�`V�V�°N���q�$*���$C#B�)�b�w�3>HL{�ǈ��gޏ�"�>�D�G��p�}@߼,�v���f|<���6��g�~Y�v�tl���JC���d���
W-�����6rH�URc���f�Ϫi'�;���FgM����R��OϾ���Q�U�DM70���-&�Ĥ_;nȹ�´r8J�e0Ŕ�s=M;;�wp���Mk̨~nsUX;�O�l�d����
Ć&1O�5����%C�T�/݁�}$0�C������߮a̓��N`�ȟ���� Xb��a����VX~\YȐ�}3����~���p�Z�Y���%AO���
��PJy� c&��Ri�y57B�S)�'�lO��>�)+
����:٢nR�EԶ��9�������UW[w����u~^�>S�<�VVI�5�U��nnJ�0*i�%��dU��X�DV���VO���?3�I��in��!{���Wu�q�����ǜ^Nmhg���LH��1�X���Q&�a�u��m�R��&$U�������*�P�+���5��:e���L�b����Y<�1����閸�_R1��d���0�ס�>����B�'�,���7����9�>��p�m�S�a��q�)�2K�f�m)Dh�#�~ �d�U�(.z{u*C���z���s(����� �ԩ'���B�m���q���'��Ъ�G����O��!���1J���ڂT�cQ����
!J(�YW�<�l��mM�-�h��w��u���ID�dd�JI�ՁX�%a+-�H0'Ԉ3���>	�US��(��bȴLy��z���$�$���$���2�6a�_��g^���kjm�,\չ��6��ɶ��iUU�,�&&�f�4=n\4�*Z�D�mn;��i�����6H�c$�>n�t��,�ĤZD�U��U�X,�$+6�6�fÛ����c�vFw�_��`<��$��v�. iy�*���1�H� �T�UQ)!�֤-�b�%N��
j��{����� l���`�G���7���WU������J:'�%r��6T�ڔ �΄������k���p���� b�F	��ݹ��-�:d������fu���.�T��L��ײ[�0�/��޲�#`�B��m�ޮ�pb?7=���t��\��7�/���6,�p�<���0S̵
"���t�������/T|v�C T6?�?&�
��w ��A[�{���<�ݓ�Y��'�S���7p*T/�(�s2~�m:�Q��l�� Ȫ��`�t��@��64)zbK���&"��A��mA[`0.ˑ¿~�)�m<J5B�;�\�좪�HK��$���=3��	b� � ynٵ�8���z�,#�����v�������0�v?��r���ӿ=���~|�4�f)?bP}�� e�����	�d}�&* ��(+�%��^������S����a]*�@D4}�4���?!}�T�q�~ b�>�AW�Lؤ ��ũiQ�q++VZ�C�_�����K��c� nJ
mtF���WH��;�ª"��0J�T�	t7�
�]���@X�aն.g
�����ܿ%�����3
����DJv�?=A��{���c&LA`ewP�j3��?�6䃀��iM?�T�?����JB�*@����u� ,���j��+B�������?��G��r� ~#R�i*�JDտښ�Hu6�NV8B�H�@A�;}k�zBw��Mot�w\�j&6H�k�e��^�#y��;]j�}|�q�`��ED'�A(8>Y�2ehy�[����A�����������5�����&��?z�N���A$U(�/��\ɐ�ȧ*�O�ŗx�߉���#��t�og*��(��!N�H|	��;���s����k����(]F�7���$d�%�r��x嵊X��`������j��HA����{�!Z�(n5'���%aw�S0����'�.��W�߻XBH�I�����ۯiUe��?5-v� ���q;�+���:�G��ꡪh��\׽��"��6���a��s�@�CI�V�v() ta|��{�<��\�G����G�r�?�)1nV�nH��=�҂F�lͦ�55��3fճkm��"�Dʫ��<��Bo������e��,S�T1*1Q�("�.R���ҋR�p���#Uv��39��ۜ�~��.�?�����%�M'U�>^]i�mmf��m���ܙh��$���p������d����)���ޖ	�D�$DF*��VDLڣ�؉Ҥt�S
b'Iʻ���$�)��WU[��@�K������)L
aUJ�s��%���善���S0j��snQ��|h�&�m��>d��Ϛy��75�ڭl]��]3�^��u5C������;-W�a�y��DHWA+��2Y���'.������L�TII Y�Q1�g8�_m��)*��UR�&U��'��.�t��XB}��I��{�B��#��E�O��9/����^J����b|ix��}��$��O�"�R��Qྋ֡�O��>��q��B�K�5Q�Gz�"����7�eE
�(1*�{룾y�ٵ���m[Vճf�~��wѼҿt��G�{"��h"�#�cH�D�d5���J0b�`"0f2���lb�b�*#
#*VDTQlm���k�UA��Z�����R�"^��3�� �+h���z�c����U㥵X��h�+�yO1�U�颯�x"(��(\ �<��_���V��~<p�"��q �562�:5T4����Q�
]��}~�$w�B�
�٦��y������3 6��������M?�TX��=�ȧ��P�sWZ�z�]�"$Wg�b<�B��\�-�U���>�=j��+�+޹|�'�SԽN/�-���g����9�p��c��#�Kئ	��Q��j+�Wn��`kbA,C(b"8
k;��
�JJJ�S__=����O^c����v���D��_!<��K���z Gex�z�'�;�ӯ*z�zoQy��D�m��t��$�IHF����z}O;�/k.kjͳ6�j�O�nӵ=�6��[�>���������{I�/������
\�0�q�Y����\����-C��	B~I���4T/KʠT. �毧����^'���7�^���E$�*q1�H������lm����.V�|ܶ�����-
�V��dR��6�5�J��J�U���ȌV�JċU��%b�ł(��
��f�Ͷ����'�כʝ�v�g�Q�:y�����t�[��-B���qC��N~I8�0a����(�*��("H�,V��4�f���E�;�sL�{=��xB�	M�΄^�Z�ª>���OW�!v�K�}�����rb��������A������=�>O���/�����!/�H��1"��ufA�^W��i�$�����A��ORR�,\¢�� d�<D�)�v��gpw�-m,�s��Sĺ�͔�J�ة���hu���'��t��iV��]Dp��xj٬V�\�� K�����8�n�\�q9/Dw.�����g�{S���5Ki0j���wi~O#�rͺA�LP��9�0�R�.MYu�z�T��A�h��`5����l����/��q��4\���f.R�m?L�	!�b�(���0F"�f͚f3Z�fkk1�"����"��!&�$��T�YtVK�m�7�k���Rɤ��;P�O�H]����R�VKS�e�.��R����tWRU�.���ǲv���]�Z�{�]*�k�.�䡨凑�<:�R)�f93^���2oЊ�
��!1� �e��	��1TDv�'�@ɢ;ʺ��#�?X�@y����'����YK�x�<�
"�U^��>_��.)s k2pL`A.Xdkߍ΢�M�Tͅвi3E�Y��)�T�4\���=���m5Y������G�u�G���X������r��������.�,���N=��ćS񎳫.�1�b@�a!$�!$Ǒ���2>:}
������G�\%�-�\��H�_&�S�UC��{��$Otyx��_H�T��.��Sx\\I��{�Z#"(���:�w"�4Cj���O��!aj8����EJ&Se�Ў������.���i	�21P0�=����]�z�Ԏ�L������x�&C'�1��z+/�v���E��E!�I>�����-��8O��Ǥ�E6�7��׌3U�|�������O��a�S��u�8��;��C��#n��%����<�<�{%v�Gmzɥ:_���uI�MW���;��v��B���ώ����"Ej$o=^_=x�D*��a�C��Sظ�2I�;z��}Y^���^�z�wC����
w�}Z����&JW��=��MR��x�sKS �H��h9�O��g�br�LC��Ϛ�|P���$>*��8�(��3QJ�ۦA�sը�&���u#�����[�'��q.e���)�������]�Fk�V�}��-�G�]-Hj��߽��G�f���P��[���P��eDr��1��/x�)�G#!Y m~�oR�<�8�K��IHH�f�9�[�}�����338F۵�
��C��;��s�}.�Љgg�w]X��)qMk8_Z��ֈ/�������\�|z^��$@!$X����_>����|%��7X�q�U���BA`�DĄd�$!|�:~�9����57 <��䄒1# ���?���� �2C���!yP�`EU"�`�Q��D]k6�r�4Q���6��o�}����h����B�����Uƭ�Zk���y%h��}�k��l�h��J��2�|��N	*Mr��D�d${����<�����j@��4�i����4Z�pI�l�c�i+?gm.vVp�8��b�vX��T��>Me�RAMߟ�z�����yp�_���jUT�l�Թ}Cp�|�����������sT�u[�;�uU7���n@��-�~v͵&�|>��v�N�������h���RA@�cK�7�y�����[_��U����K�{��2?�0!HO��wկ�}�E���?��	��յ.{����އ�� z�7���&�)���%��p._p�>�h���wpݸ�ǯ��d�Jl��ﶴ���bb�x開�V���zo��h5]��ݙ|��v{�ݪ��_�g����7��7���y}&����g�_��%KX�$��4!k������|O�R�����gn�]����������k5���� ZDH�)�'�9�RI��s���!lPY=P��jG��4�b��N������p������vΧh��c����b[�jv���x.��;���������;�UsQ���^5�E1�o1���t��HP���<���R�Տ��q;?�w�K��vn�k�o��u�u��>떯z�rw��y��߾���Y����?��������~������ߣ�^����۵������>�o�}�0��}���������u�����[�W�?��zߦ��Q�wSǳQj���}�pS���D$�v���?�y�S�z_�^O۪��o�=�������
Iߛ���C�Q�M��w�q���M�D���|o�T���*G_���_3g��}?�_�<e�G��ϯ�~_��\]��w��$Й�����U�ϛ��Z�?����|����d��}�V_��U俖�=W��sYmk��>�uּO'x��%P�8���~�2Fc��_�����3���7�Ƙ=T�b�0�r۫�W���,��S�OΟ�~C��B��
�����HH����&�o�@���Y$a�/��g��F_ڼ~�������{��x�g�w��?���:���?�z�V����o��e��߹�p}��=�_G�7���J6�����(�̔fŏ���ު�r�~���O��B�_�2�~H�pR�H�#M9w��X��=�0��?���o�_�!$���q�/���(��0x�z��I��o'��>g��_O��WM����|�.��Soʯ�O������n��u�/����<����6Ї��S�\H������?�$�_���~��3�,��P�o���o�?v�����g���!~r�/���[�\��f��/2G�8B{?� Ps��i������~#�k�j�J���OO�e�؈�/��?��s�!�����I�^`o�j@��8�	�"������>�@w�C���v��X��#�K�L��l]�j57�۪�F���jD��y�lބ��.��s,fH��>��>����$��a�����9��0^5��ƳUW	?N�L���I�zO(֭'Ԫf9=�c,l�7
���?�.��1��N3�=
��Z�.~̀�V�S���r�w�˳1�^�	C���A^�����7��`�[�=J��d]��L��$8w��y�`f��<<R��A��c���ر��v��ki�C�T��p��(���9�nL��E�b����m���z}!��"���B���|�m &���w(o�L��@�:�/� >�T'��*\EyW��9�~����YQ:˅��YW�U�?�i�5�O�g���~z;��.b���(�d �3Pe��B\�$O��i���_��/�?o�?���������?�����_�28�+���?'���}~��'���{�'��<�pv��I3��Q�;<?���;�N�W����S;�_�a��e��I?�YP~���n�2���q/��iO�#�,�����>��?����=��������V^���4��_�ֿ��������?�_�}���7�>�����>����w�,�������A�H	�fx ���:�����Oճ��M�U��J�q��F�r�,#���I!��0�[y�/9����_��t�P���̚b(;�¹�!�M��J� �ӇR��Qbe)��sWe��,�w7n���i��f�U�~p}���Uo�~���~���}��_����zX������������%��#�JAQ���T~��Y�����&��ދ^�CH��ȣ�㻢�:��Y�!�2d���PI�_�)]�w���a���4���^'�v����d�M����;������w#����M���>���0�'�E�&bV�r�����i�����m��x<���q(�����0����!�4F6�D�I����g:�tFEl���ZHSQȝ�O��2f�U7��  �����SA'a)����M��A��ۧ
�� �ޣ����/vv��td���0��c55�YI		(����\���c���V-ojڹ��S��ӣV��:�1#�2#c'��?��0�� ��/����?���-(�����b"��U�Xd�W�3i�p�d[ 2 H�yk����������?_��;�$�b��'G�y�(��,�����='5�����[gԳh���'�뺞';�k��W�-S�|����o��?/c;����b���*����r�
�������������8���h���������z���D_��Z�?���?���?���W����~��~�?'�0}���䷔q���M�7��#��������	��u)���������͍w﨟�Փ�]��̟+�=��������W��56�	�U��"��GY�ߣ��q�����ƿ���'��2?d�ُ+c��-�p��HE�da� ��Nɨ�=M������Gڽw���{߱w������a�����\~Ez헱��8e��R���H��v�����7� Z  #��� �!Qٶp�~霝.�,�͛n5�}�����I�K�Ħ]h ���g���@nEEz��B�R�MFKj?���2��I�W=���V�և��m�}.v�����l�������+�l�B dXֵ��b|od�;U��`��O�fI"�?��,;�l�I& N�];�ٹ�G���r蜇Vr�B�D�&��\=MdCn8?�|��mK�Iy=��j�'���Y��8J��%ՔK�TdA��}��&�����أ�"�`���o�<B��Ac��+�8�Ǉ�v>���x�����d{|�=w��},?������X�ҹ��o���G����3�{^���\�o��uN�b���6�9����\VG����^���b*�/������z���������8�����|����~�A�"�֜��$OY��c������� ��*�(�a��S$?�Y�o�����D�zMy�_T� 6A/�<���@�� )��0{��-��޷�zn2BZ� ��~���+���ިP�w&�P�T$�w��:���Ϛh�.�O���,�c`A�Ȩ���{����5�_�jM1��6�չ#�J��%N쑰���;NX����:��?yD�7��5���U��� r�ߞ�*K�}�?�x^S�ڗ"vۮD7-��P��Srko�O'���~�I:��?n����Gm�-j
ؿ����jk�*�#�~H~��X�9G����c��ǲT��_��Y� !�w��
��ǯ�F��,-�����񬲝��|����vsbэ��!�v��V��j���߹�Q��(�Șp�m�T1�_˸�*�~��9A���j��ij���sà֒~1�O�[v�U6�����.�D�h����nWUcKQ�CT�`�hd�A���W���>��w�m�V��9�ѩU�Dd B�}H/�Κ)kt3 ��?s�o���߁w�3KQ�eZ--S+I���`Ab*H���6�����/�o ^b H	��!D"#"#ֵ_��!����d#	vG��m*�E����C���D�D������gk�SbԵ0�be2�10i4add�7�t��bqN����~�����r�h��y1O$���M���BP�%(R�4���)JP�]�)�?�� ā'��?���Wn��.�G;���x��ܩ��0ν1��i�|�;�������E�{6yݚ�����������P��S�� �F"$ �%�_�ET��j$�)f&%���o�1#-]Ю�h��V�˫$�w"U�2��唍f_��W&�^�t�G$`Ԍ��p������xR��j�:yO��BIi��UY��H-����Y-F��+S#)���>���XAH*��P�U�qZ�0�c��H*����};!}3����|�����*���wj3�twؒř�����C��B�}>�G/�r~��ӱ�\�h���S{S�}ny3�t.�����q���v���-/Q^�� �1�{�e� >������  �"B 	��&��:k1���C��Cm�J-�bG�b�	�b�\f����2���:G��Nl{�e�l�EL�')�\"*S�����8M����-{&a�%�+(s�k��g� ׵ �`�+Ar�R(
B��hJ�4,�d����A�d���:=�Z�uJV1�9����=�f��)U+R��!Sy��=��1�a~�U�~��u�m�L��������̚( @  ! ����k㐁�x\11Ĥ��ckX��8��bWzҧ�H|#��=
��ing�ע/�ǧ��TԷ��33o�ou�dA�Q`*�c�X:w����9Rn|��L�����a'J���O}�C�	�]tNB���:DkmƽVM�И�'�QrSt��q�v� �&)M!��!`�y����h�CWB�z�c>�)؇ܖ X%E�I`��-���JxN�H�s`�R�.:�G!���bbK�;n��*�!*��   3�D�cj	*0a�����]�����#���k����̷��n�SZ*�DB;mC.��e<:��+��a�s�����^� �8��Q������8�R0"�7;�,�7�$x�}���B��
�V��M4��U6��,�y_��۠�oc�`�NP@g!�"Z�"�0��W��e`�KH0����tE���pE�K�!�Ԕr���F��Թ�䵮�q�$��)���Mcy�!�k�8�E�V��g\�d�u�WYB�	�x�9��l�V��9��@��c,B� ��)��1$�[�vc�<xb"![��P�7�����erHʠ�E1Ab���"�ADQ"����b±ZZ�E�c"���,dPDb��fM�m�ҝ��M-+SQ���j�m� @�@����}��@Yb��J���<�$�u�H�݃�����	-E���~���+o���5��U�ՙ������E1�X��K�j)Xi91u�T�vx��_��p�Ko�Ox%��i��垺�cd�+�3����N6���2�ʹ)��V.�P��� 3j�:J(q�>�9�r�Z�Cyk��E��A�6:f�ۜ��%�N��9���V�۹R��I���ޫ������L��[��5V1�P�*��zl��S��o���8吶1�%�4:����6MĨ��3|��b�㊯x�ɹ�R��]����,��=m8/Z��f��U��@*/���-���Bm�����N�m���عṵ�a��a����� � 8 ��H �f��G�V�B�
za��\V�
��ȩ�?��n0�9Om��Z=8����KX<��Y����ꮐ�+v���:������֛kF�\��Q��N{e��\��l1�f	�%�,�~�S$�T=K
i�p+.�h����1)4�a�vrZ�۔�[is�#x��� 83����80�[�ң��W,��Kva����\t⌊?0^Eh�iF�����σ�
���x.��1�r�++�[g�NWr�~��%{/͊�\83��(%�0�5Ti�r��\�f���Si�����m��ĵ�a����d�&쟟\��S������_su��x��C	���i�@�)`���d+u�p9d��`��e��כ�v�t0�<��f�-�{������=�>x�p!?��'J���@D,����
�e������W1���ת��r��(��ÏA����l}�3�����
kp͂*Ϛ/�@�]�x�[;�[��)�r�B�����(����Im;�S���ax��֥m�~�{!fNt�ki��e�,�SU��<v)�W�7N�w<��=�>#��H�tx�B����v.;�ӵ��M�^��+-.�ʳ�p��'R'��wc#�l�:�a�أ*�Sۺ�J�])�6)��Z̶0_x�a�n�7-�,L]Ǎ��v�|2V9�>qR��4�uʣr)s�4F�nW�r���������[���y񽵳���B�"�-5�vV�]���0�}a�Eս��n�诹ie>��*(/E�-�����J��M����[Æ�El6�˶��;���M2�Q�;=��(�p����hvF�H��1�g+��l1on�M�ٷ]�4XeIZ�f��j��ս�k��5~��월�m�xGH��N��N ����� @  	�   V7�q�^�[rJ}]?����<���B��>�=�ا�S�j쏉ӧ=`��*[��R��Dn�Y��[,�|Z��)z<3��^�>O�67�����ek���W�FC\:�9��8�8qJv~2�!kygo����������f�1V�|f��7�:��E�IķA�IM�9� )h`�Qؠ��mz�oZ�����疧��޽4�
�ߵn8w���U�z$���U�}�).��e�j#��泃��7��];�۪{v�r�H&�Wa�V)�~�xy+�e���'���CR�,ܩn��V�a� o�)��:ۻ�l��xxe�Z^������wE7qY���l�~=0�W�w�½C��g�ۮ?}�:i0�7h1�8Ų��y�{�����s�:�|��]Vܼ9n>\t^q7U)�kpӂܻ�k�]�S�&�-�[��^��n�zwh�S�]�{���iH&f=�^&�yKR����A��[ lϖ�qdQY{x�{��0� 4!�- 	��E��Ҳ4�V��)���d�j��^  ��4M��
c"��u`m�\����
�X�@�Y$"\1ms�@�^�(��6��A͗k`���	+�l1��1�"��r��iRG�q'�Q���.Pa��� �H�=<�K:�
ѭA��+ Hh�!�$ciVKlu�-�QUZ-�'f�W��Rf8�D(���%:�YPȴ$8$6�	;��,�������\���El���(yg~���o�^�� ���+qZ�&LDZ�R�0S|���	��A�?�Вӎ0��	�J��QJ��}�+9� UiJ�]��B����FJ�,�*����@��T�)T�'x� X̼� l���
�N4]l�����շF��c�ޕQ�����eݍ�+��-�ӭ�X�Z���Hs�W���2P�|q*]�yלQ)R8�ƞ�A�y+VgW��CM�I������.p�4�j��&�=�"۬Ue�m7V:ȕ
aO��m��HM[c�Y,�,��d���R�6�E�D�7�J킘��Wt7P���];��W�۲f��c�R;�G�֒��y�=2E�e�x�*x7%���G;����ƚF�ꈱ"(H� �  x?u�P+"Gh���g�UE�h�}��x	��J*?�qa�z]���U3M3�	tPo
ץ�8��̡nrtn3��V!�6q}�x�3@)L���$&�E��P(m�V>��9$���P4�g���j��PB�F��FQ�v�td&V碭
�Y�!VԑP5;Vm}��fD���\���]��m!8hj"Z�O �(� �<D�FBO�^�A��U���o\���漇��a�R���s�# �xc���ž��S�B�R9՘��k6ĸ�L@�H��̅�6�a1��(|����hHP�n\�cgEt!�R��Y7E��D���z�d�H+L�1���`4��bp�P��"i���.O�D�L��+��&(�1%G�@�ؑ�(���<C>!��`4y��P�@2\t�c���ЦZc�F��n:xM�C�~W���pB���e�p�=�#�p��t�]>�wS�;IC�̐��4�&�2t��(̉;�N1@YH2c�`d�%��#i2��(�F��uIL��PO*�w�X�8�j*,tW���0H�Th-"C�\�3i�>��AR�;`]�����Y>1�E	���V@&�o;%f�r��Ln~��ڍ��o�o[���򶙦$ �I�I����@hdD�RDaOY�h2��{`�IU��`�2��:�:�$ hg�@{i��M����-_]YFD9c�0%kV��+0E+����M��.�*8�AXa=���o8{1�����/S4�� >}��ݤ�`B!E*[ ����\E�Ȇ����s`�a�)P�tk�j�G�|�qb��ۣ�pJ�O�qO@��F�p/�hr!�n%�� �7�*'0Rڱ���m6ѣ�2��,Oy
}���Zژ|�Z4����+�� ��\�̪I �0(�f/�\G1�E��w(�D��4`J�"�3�k��+*
T���P��L�M$��������<�P�T!A�4��u�\�l�B�:ڦ=�6�8�\�@	�h*�%�`me�v�(�`�Q.Rbj� ;��7Um��0�~k-tmuSWo*Օ-\0���K6^P�|&ݮx�����c1��rX����dI=iE`���쨊I�rf���(�bJ��5&���L*Vm`:�)�+�tKӢ�� 1,�έ*�wB���[9d~r$rMl"֙�o/`�SlK
�EtTiIטX$e�0=���~9H]�"f�e�B4����ڴ�AU�2��d]q���p٬�W��M^a�c�0%�'
��VJ$#vi3y��@9p�۠�f(��m�k�ӭ�XEL��M�U�g���&�Cn�sXЃD�$��s]� C�Neq��ߗg��κ��5�m��YZ�&ΪeI6�N���t�8���AT�YR�RYIjHe@XX
ň��B�kM�3�mm[\�ml��[+i�m�!l���E����TF�Il���Vʊ�ҍ���(+X+!Q-��A)�ڶ%�M���0��H�TE��-��S13���n�ik-j�bfT�r˙�R�*,�HJ�
������[Q�Nd�sC��dQTX�RE��TR1X�,���1E��d�T
@+Y�))�)Fռ�ŵ��mVØh�I$�H�Ȭ�Ⱦ���8?��y���ټw����~�~����~����������*ϻ��G�?��O��u��ߓ����\ָ�?���+�|����}��r^6����~���j߮z�;'���|��~g��|�Ӎ��oA��^����\��|N�n�¨	��F#��Ȍ�A`�
,EdX��b�f��V��ce6!���6KjmCV6�e���ɚ�6՘lڛkd6��&ͅ�l�6ڦ��M�[M�e��Q&��)�A�b�m��-�D�6+4��fڛ66-�V�[6CciA�b�`�i��l)��cf�fl�cm���i0��TTPEDX�1Xkm�6�[Fɰ������6h[�M��6��-�lU*��m�l)����CbmTض��6�6��Ckcil�ک6fɲSm��F��M�M�lF�[A�6��U[(ڔml-�l��-���-�ؖԍ��#iU����j�[&�l�mҭ�mM�l�d���6�Tl����UmJ��hST�ڇ�i%�*F��4
�jUV���z�g��w/k���O��S��~#�~.���_����y������_��o�]�0��/�w�>w�?B���?��������Ɔ|���?��� O�t^���M���>G��z?��=7A�q~/�ַ?��h?/��o_���7�t�w��q���S������zڿ��ܯi���������?d��v��~?C��Ӻ�w���-��������7�����~/����G��{M��o�k��|��u�����3��{�w���T�]�o��<�C�x��k����$i~y��A\���v4cD�YB#(�b����QAUUVEUc*1AV"*��"��TE��EQX�A�(�EQQ*�AE��"��DQUb��+
(� ��2,dQ"
�V$E���"E�#TD�����EQUQ�""�QDATQ�Ȉ�Q��e�mZ�c4���X�
�dX��H��dX"$TT���b�b�*����bV*�UE�TPX(�PEAX����*1����QT�Qb�"��PTH�UAD`��1,U#�őb,A��E��
"����� �"��
0Q�A��"�(�UV"�E��(��Q��"�`�QET`��`�`�
�A�0EV"�
��A��F(���("� ���Q`�F
,V,QFEcb�U@UQ�UDV+"*ETE�+�
�EX��TEb�����*1P""**1X�QQUEE��`�ETQE�+E��TE�V1b�1D`���(�0A�(�X(�V
Ĉ��F*��#$!	�����J�|o���Z�c���?'���7��V�/υ{��=�f�wm�-��S���_����/X�7��u��������繯���%�o�����N���>���=���>o��������w�����ET]�R�

@�H!�����;��e�����]�������j�O��p>)�����y���?~��m\���������~�o��~�|�~~������W�c�����u��1�".���>ug���N�~�ϗ��Vn�J|Lwڻ���_��^��buX�ݻ���J�+���}���g����4W�J;°�߬����ON��g���ҊB ����x�"	��0J���<[�ǨVS�6T�/�=��Di�<E�k�h�bw�Z��Z� e9(s�T��ؑ6	�~�?��G�?	�b��q����b��o6�c/�+������{P�U�xOQ�S(=Ä��^�-�ɒ-zI��Nܽܲ�a��̩��s|k�e�t�e9�qz'�i�j�E�NN�`H\�8�B����$�:���Y,x���s�@�\SR��ww&��-HcT�!MH�	C���LyΛ��됛�F�q{\lKl�:��?s�c�'��	��1L�U=��`8z1$��0(%�U�1�S�>󼁴%%Ya�r-�M�j|���4���w�뭸�3�p!j��!�X�����VBe�j|�È�JYQ S�#��-i�C-O?CWq��VR�xRv��"�7pl��Z�z��qא=��(��������@��sIq���VŲ$���T3@��v����d����G� wiV�
kk���l�XʨU��ȬIC��aB��o"��:eIs�Dr���b��B/���A�Y&�Hi�K�ܛo"�G>+">`5|Qt!A����ǡc���0��{�n(ߩ�p8��^n$��)��:�+s�i�cJ���1x�c���~ 0/���L$�؉��� ��h������_g���s~�)θmV��:��7kg����<§�����w�Cɉ���1�l�a���Y��>��g3�YY%|�a����O��S�$�HP?ȸ��k'�Z�C�>ЁY>�d��ό&�XV�J��Hk\IȤ�����EV|d���VT2�=���𘾘>V�����U1R�r���+��>}��P1�>�7,��e@�{)1'!?	7��A@��%~��}0�	�/& [�1�?v��=�Mf�_?}�ֳɉ�!�(b�`y "i���18d��|C�dĄ��O$���� E]j��l)v�v�&�A�\ԡ�#����ҁ��)�(��A+��Jl��l�V9�G0�sNeI���A�#����֝e!�����%��RWY@��^8�^�-��v�6��qv$��/E,�� a¨�"�$ߔ��d5'��V��b�>���~�y>��'���É`C��PY{p��^k��g��H}���`|B
C�I�S� |d�"�Ր�$�1��P� rMO���9!�$�B�����<ȲI��9��2�!��I���ʒL�[S�x������v�jy2��ɻ�m\�᧭=J����#�9m��[6�lڶ������)����ÁJ�������������������������������������B�&ʐ�$  E�*�+�}��{wN��=:i�mF���8����v�=�@�PRR��O��HK`@     x�]�����}���u��8v�Ǹ�g}���������L������u��n븨�s5am����}����2{ݼ����g� Oe ��]�����=2�lkY�w}�
� ��:   ��*�{xz���.���\�;s^^�n�WP���:�{r�GmJ������f�y��r��r%F��e"��Uk)v1�ݻﵐժk�����,�kץG5��z��:����u�kW[�K��S��ngz{#��v�v��
��  (>�   �m:=��q�=��׽���zb�n�{P�ּr��-G���=���}��v�٦� ڹ��^�o{g�h�v��@���>�!�T4��!�=揻U�ϗ��%'  ���gɛ�����[0Ow{�����ovN����n�{�����\��3n Ç�O���h���4#���y��v�o �<;���w�G��^���� ��OSt�|          ۼ 7޶wwPG��s޻vy��{���������vڀPTR�! 
�R�����S��-���"�Ʋ���n�wu:�lF�E���8��s��:�+����t��{{��;wmt����u�❭�Y�i-/]�K��ͱ�P���nݫny�8�;��;��dVَܜ����̘���l��I��m���lƨ�����ڱ�� ���":�f�+n���ݹ�բ�T�ڻ�;
:�kch�'r۳bMn�m��.�W�s^�t\��)vٙm����U���kn�u�j��׫ݻ�n�,�r�6۵���]"W�m�m��mr�+[����W�v�]�mT�m�־�f}��,����s��bz�{ۄ�����{�Nx{�B���A�m�h�&@  `  &M�`�4� �M I��cA0�L����� jyA�  �  M 	�4i16�LF��ț@i6#Md�2y0�i��L�ML�h&�� �	��	���M(� ���h�CC�d��F&S���?QM�&��$�j�CF�Ḍ�4=L�	�z#�����4��=4��Ѡ��Q�4?T�=@�h�H�	�@ �F��eO�F�3Q��4G��104Ҟi#��O�  �3i��4zM1S �zh�4�z�A����L�z�$�R6���4 �" � LBz@�2 i<ML12�D�D��	�&m@�F�����*~m��cD�jx)�S=��=4�z��=OT����5<j�ҠD��L&�	�&F� M10D�di�3M���(�4j`#L�a�=4�<M�S	�m&��2M�MOɴSɴ�C��E<'�� �$<�� ��Io`㒋��D���ulQg�&uy�?��~�{� ���2j2�3�#af�>�M�2t�`�0f`��v�նv83�g�+EL���H�l�1����Z�Aj�����o=jҖ^r X+C˺��e���Y�k����#:��B^�������Z��F�NJS�q���g�lw�qdR�2�V����+�T��rЈھ�����A��K�d�+ z��t����G�����c�[�����Q��>��Y���K/7�X}
�J6��ʵ^`OHx��;�Q�����\y�q�&!�3ؔp��fX͊��>��{o"���/��0�匀^7�)�Z���볦�n�Н>�3��}_�����<�t����3�3��/����K�=�zQ��Q�]ن�������}�_|/�6�0�?X!;;@��Nъ��m.�M7y�}�X~p�x���a�@q�;��}λ� �gӡ�6  z"͙ҍP/U)
���Q\}��̐.,Ѭ�7e!���ĩ0Cs̕����B�ê�3��Hh�͚��kkk�J�0��0S��g����I�=�B��J,�]Sl���`Ѓ0����g���B���%�}�����a�X��e ��B����8����F��2�@��<�؎��O�r�՛��6�H�H�v3��._��i���������*iAڿS��OoMC����	��彎�A�V��Yc��w�w��yǖ4�qH�M�l�ʛoa_��K����{�@�L	~��V�/W��U�n�����:��:��W��o��;��]0�໼'��9�{��P��/1��
�����co��=ďHlF�QMe�X�m-t��o$WL�"�p)��t�]	i�!-���܉�u4��֡�%,���O�D49�W�_Y�P����p%�(X��2��kWk�vg�mx�\�á�2fm�.�4����!�����:t�d��o�WU�����%_o����ms}����vw{:�����?�{�Wfʯ_ö��7��;JC��I�������^��&D���9�K��x��)��L�/w��?w2C�[�Dwr�{�ĜŅS؇��Q#7��{3�{Nu�=)����=g���<�V/���i���;��6�2��EȒD;ħ񹿇]>Y�~�zt����A��Owl��`ޞ%�����9c��^�t��/�����x��@��jGA��γ�z�_���Sק`�T����e�Ni�L�:l��>p�_M��#2���#�k-��O�:p6n>)�u@���5�}-���y�\,�Vu,T������$ߐz���J����{NZ��]�����i���S��J]C���3��~��Cۏ�$!���r}���"/���E ����lг=b^�~��$c��oF<	ӡ3��&;O���7Ao��Ȕ�����Cϼ�v��וPE���m2Qr=��ʎ[���� u�1�C�D҃=��i�;ܽ�A�(��
K��h�|���kןk�&H��!v�t�?���y�y^=��|]H����tX�3 w?x-aŧK]�
�?��g_�]=���|�>�������]�c�>��S�独����\�>�Ǹ�|�u-������̎�L�;�#�ϥؐa�����>J��vk׺�?�:z7�I���WW�'��Yzļt�(�(0�N���"����GK�I�q����õ��Q����CY�p��'#Ei�Q9��u�%�1�
��~^�>�����kt=��m��xEú��>/\��!t.��S��p�m�?���}�����:I���<�O��������.;:?�.vE۸��wA�=��7��z��p�>��y�ȻW�;z�ԯ���	uۡ��ѥt����CPN�c6�T� I}S��XT�'n&ck��\.���)�DKr�SI����3�⬬u���y(8����B��):�zFȁ!j����S׊:�7�����7�@��uE��=��}����{�JQ���K, ~+����*Ӭ��]�y)nJr���>�I�eF�H{<J��~� w���°Et`^>َ�0��-Eh�A[c������(m�s(Zc"	R�����^tP-;�%�]&�F"�D!�e !f؛���<}E�=�u�Ku2-���wO���^7�Mߥ�#�ً��Z��/����Xw�+� "}�@��/+�rlV)�-�w`�KΓB�؉ϰ"b�q}l�� �K����Z���̮)C�o�B�C}�5�Ao�d<�_����:�{���
���k�?I񻋰X_������(=�1:��dN��U���XL�1�,Սs�k�o&D9W}Mt^��I�c�H�hK������o.�O%r!b��!^���j����P]�M��=�����raW2��(���:��מt��-���wU#уw�^�����ؿ�~D(xG�?�K��aO�?E)��|��s�<(��>�n����zW��\Ն������l[��<�9ZP�J�X����4��AiTk�\�XF���b&�};v��F�Q00�Ɖ�&x�)���������iGCrAXG�tx=3�n��� �p��k�$�qt���1�Ñ��T����cJ���k"s�;�	��>�E#ң�����Y`ﾷ]@ł!ڨ�.!�[��S!!��j���5�^�;����]E��3]f����m�sk�yCm�c ��`�I�����64��[�1oF�{���A�g��7z�O]lG�Pv���X{J|ŊUGHb�ު���oKY��1h}vd5u4��X�I����~F_�����=����������SRc�����n{�مC �-=�q(�����N��g��j޻c'Â�X�F��A��ϊû��2`DN��;��2�!�t<>�|8����с�0IUlgg������h����0��Kt�ұ,��<�LPWc���wC�<{�����`ěZ}m'��_�+��E$	�ncWtSmM�pSΩ��L�*hȦ�B�e9��1�"	�L�̦*b���3'PdTb+ �����NϢ�p���棖,"x8��B�d!@X�ګd#,�3S��Z���\�����2�ݪ'��X�T�����1���f*�	��5T܆lu��_ޡ�J��J�"�q�e0E'��ܟfw|�N�DATUATUQAda���5���!^�@.�eK�D�³C'G��^I����8���*�a�9H-v��7w�����'�ǩU��f�Y�X���le�g�n���`�8sUkW������������l�2��1��I6D7�������Ow�P��������m�E��PS�R�"�߲ye� S��y��~��fn�T�Q�$z���G�B�ހ���=�S5������YL��	�% O	ʲj�Å���#����_	"ZHTf�ʖ�p+i(��k]tڦ��Sߘ�i��S������)��漎:��^��d��ܱe��w���ބ/ȣ/��͛�6=}�� �����R���R��b����_�X)��iJQ�$�^�f��u ֢��8�mpÑ��{�/Q��pu&���Jh�s�zl���f�ޭ&�T�R���ǎ:�&���i��I���QM%7�{�3^���(��u�խ
g_�Gߺ?�����kT<��cg?�.��nj)�N�|�\�ٮ+�ۣ�w��TЦ��)����ɧNC#�8��c�G����?a��S�fCM^6��]\��4��������϶\�¦>��]��(�,ë0�H�� �@?������e6Ԗ����X��׬�Opt�2�Ե�M6��,q�'�۩��� �_���=~�:�o�ò�p����n|���W:�E;39p��QN{Z3��@����Xl|�x;寸��0��d��1���7M_���pێ��ax�A���v���@A|�D	���&�Q���\�������طSƳh�[��B���S�Q`�z��Am�%����/g��ύ$��F�oE�v�WG��q����~�}_@�f����Z�9���ۘϊ�|g3��ڮ��� -b
d��8�yl�&]�'�ۯ�(�PQ�E:ji�<S�$�SJrjܤ;\�6(��^�ćk0ߚ�����p�*H���;v�cN�&�b�Z�'�m�6�d��IFh��K����c�.a�Y{���yk^�6�W�U��-��V l�ʉ徵�����(����
j].{Nc�����d������zlm��2��lY�Hь�Yk����+����/%�ǫ��akρ6�S���X��:3�[�
��\�綶7��Y���C�L�Jh�R�����^Pv��D&~w���kiŅ跢���C�p�Ν�/LԪ�D&���c|-T���j� ;�����dO͈W����Oi�x�a�"8���{�aD��lZ�]���d�b�J�Ka���є�Fd��)�J��FaC�Lݩ�`�a&��X,��<�pn1y�M����o�%����a�N�1ɂt��t��c�k<�_n��l9�0݁^��f��;� 0A*`�A�e�(,_ջ���lZ;�Υ>��o���+Yknl�}�����iַ��01�
K�\����o��f��7��[( �;���%~+�N����8����i�{�Zt8�U��˲L1���0�̪z����_�����b ��e����:�,�mʦ=��Ӄ�[I�7�i��;�G�\]����5q��R�f���[إ���b��:�\u��R�|���������Eꚯ2����!	Dp�2�\G������;;�Ƀ�d���)���~�Rvv�ޡ�4����0��_~�����(��__7��x�!���AjN�0e���Y�l�M"�ZS�P��y�u��̉�\�*û������� V���=vI�0��#Ƅ���_ݙ0��a���D\� �,��0��C:�
��tL��|�'�Og�~uh�}�B%��'WJk4�-2�.��~o�G�t�����̛0"�m�����ӗ���_�f|ۯ���J�!�
T���\�SWe��2g5���)���N4ʔ����8��\���n3ʚ�M��Z�<�σ]g�C��]/o���@�ꂀ�����|��|@!�]���c����v��g�b���~�Men�e��mo��`�f��w|_'�^��������.�����Q�u7������ba]!�,jV<+�L�����  � $��Wah��2¶e9v�S^̍���^��Y�f�?q2�.���P�ލ?����~}y{�+۵h>�K+`"$^��z�J
����f�i�q2y�%(Ro�)K�ߙt���s��=��k�p@ O��h�L��=��*#��<�kMI,)x���7�+�;�v³=�zfB�4�Qɢ���8g��?~�f�YA��� ����x���<��9���?���/��$8CɭZ%�R0�df֮�y�l�ϥW!�ޑ2)O;���]���M�[�<�96q9�{	�՜ܸ�ocԳb��k7q{+�����_��;�^`2����, \аuIS�

Z����sRq�_k��9_�ց��V�,I��E
̥��o/���#_4t��TF�����*����2^�fEZb��}��/B�α9�5��ɣ[���w��6�^h!$�%��S,���D7,�C�j%�!v[�6=�OAu02���G�Y���h��u=溩�X�߲�$=���楶'�ȇ�违��������O�}OW��b[�`����qkV�x�6���5byL��Y�Zk$eR8��� �U���A��B�%��kǒ|K8�`�����4���Gc%�m~���f7��n˻��T�f��r*�P��+����	�h0�**�u���D��[����doVO՛ÿ���ܦ�ޞ������L�Ҡ��4 �2$�2��H��o'�s�e�9�c��A��O3���E��2�����?`���S�Хc��IJ�^�^r����SP�vC܊��dvK�%�D	d �V q�B���p�~'���-�����8gY�UO��_3Ki�^���x����{չ�w�묧��-�0��������W�8�m0�oӣ;x��k.����6a��B�?%w���;Q���ba�KO�����V�nW�@�y���[�^��^��^���}����n|>�����v��,�Y؁&�H{C@��һf���0�,FH@I�7�9����X�����]��Z9sr��O��
��.b�\��kP�\	��a���B�lR:�9�>{�������m'1h�躇����������&�� "F��a��:�!�a5��'�{UzS�u����yd�-h��:�#�w��j�f���UX�}�gJ1a��G즖��}c@ ́.d	����Ūrcy��_.ne�sg;��
~W�����F�+o����꽜��t��1��ו&�ra~�0?(욐�2��аB�>�˕.����f�K�^]��f����K"�Y����}��vۭN�!��ˈ^�vk�y������w7T�M>�[��8���@`�dXІ@�J���߻�h��N�J��1�A=���H�[��S^��S�!x��3��01`�z�c�H�u�[kkN���e/ɞ0�VH;[(G�;���n�3�L���z8�c��/����M�~c"�x~zL���e�-���L�y�۵�@�j4�@"ŇʘY������a����\�I֍wؘ�(hQ�3�<,�F` z� �-t8!ݯ�ܒ�vZ���7����/e�'�[�������ET��8�R�����
~K������(�C������"�y��y�,�^�6}G�ڴ'���my�׊կm���t�..��l��b�a7��>P�������ۛ͞<�3��>O{� ��~����2cwYb�����W� �+0 �ꌆCĻ=��v��4�Fcw����ռ��O���?ｋE^fws+_���㭆��mA������`�'��̳����DyS���߆���2c�ک�'ap� �&�L�������r��:˞�UMC����r��w%۵���L�,�ʺ1���b�q�A ��O����^��Q����t�"U�Iʷ�����W���v�wVk�?���ۄp+���W�=ͻ�������g44l���{����� �ܽO'b����_�Fa"�!���'i��A�����nF�'�;t��v��fk������Vk�'��Z�ogE���UC
H�(�͌;�K��0H�}�����>@7���t#��L��&<�Xs�g��4��CX�@Zw��c�-���d���p[�G������yQAr�,�aV`�%��Gs�4Ek���[2㴀�{N5̘�n�x��z�֏���D=\�ݐK�'II*��L>Ro[Ix���ܒ������'�/FBN�}���T�ש{jt��m�/l�\+�����8�u���\}�1�mwz�K3�=E�=�����31"2>����0���8��q-�"�Ư�т �j��29w\�_ �xL�r��_`0��Zl@u�<˽�; ������V��Y�f������آlæ�a^~f<������Q�<eN�[����.�3��z8�<ͨ�|����P@�P�A��  �0D5KIw��l=�&��|�������t 8zo�ثaDƵ���hH;F�J��ߗ�2nsq������rj��×����)8,Ǐ�`�� ������ktH_����e��C�[���D�\�]//�z���9�t��qx��#�E��?��,~5p���<�=;y� C+y���a�*zK1:w�`�p�g'L��)�~�H��s%� ,dh�6�i[�5���۸F����*{�k��Z2v�'����k4=m��Ƞ�è@�2fd�^*�!1�(f2�e^f!�>_U����Nr�;J/q���R���7�����w����H��s�{�0�����9J9{�.�:)&���eq���j�� Az_8��!�%\pX达8������U�=^XF9aSs���.�Ifn+��� �2�b�����_V�o1��i���:s��z�7Խw������4��'������` ����-z@Rf��WH�M�fr���m��q��3*;�$\���毒as���6��2�"dehb�~B�S'x}R��# ����k��D�r��~S��!-���� 0s�&H>�tlؿ�c��½=ͰD@������-�d���L�2!��p�7��g��<�D��4��SҼ��X�1��EΗ��E�c��C&"/�ųx�<}S���,`�t�S�F׵\�ə�! ������X��ў�����컭����t|{�ʩ��D�Z��Ur���-�+��mx'3 ](کEe��:PW@=+k�7 Q�ˑ	7T�!{!��h�
0B�+���ǭ�mu�N�wU,�	R}Zj�k��?pt����di.�NN�AC4��pɍ���TQ���v���j�o�j�;;�B��5�� �\d 3"`���A]�f��x�KeB�O�4�b)+�26+�,��q���~XW���ܥ�����W��C�r�H�bA�/�%K�Xȍ5�h�;��1��{��q�W��4��=R�.�OC���6��w[2E���ǋ~o�:|����]�L[@�-m�{r54�-�F����R��<W�_}���Z��m��몍�C��>�,]q7����K��{�L������_�z2��z���-W���@� ���x��G
�댚�9"����9�7V��������Uݥ��.��b���V[q��\��|8��� 3" tI��O�-U���7�\����� ���f�y���B�0��yj��݄S�ڈ�]�V8d{��Td7����;T[������a���ޠ�	X!-	�;����n���2��?�l=G��>��X�AU�\�vQ�t��� :#,�.\;�εȣ�=�������bj�����lz+v�k������x���D����1%>�T1y�����8�Ͼ�ɢh��{���9{�皯���P�Omٻ���X�� �!Z� ZF� 1�;�/���zS�ƭ�g��oN�vT.d�{�j��
�"M
���ҙ}�|k��p�t���Uq����̰v9��/�[>�(�� P+�6�;����=Ϣ7��O�/+���Қ��3Z6yP.��ͳ�z[�0F@��RԼH��趤��w|}����~����/�� t1�_uP��d���tyN�U`�H�-���A&K�RP��F` �9=�oA��k�qh��h�l��Z�AwaG,����F�z?1���t@�s�l��&��m ��.�(�'����㴂�^;r�׷�t��wZ�a�{���G3 
��_��a��tq[>�R�n��(�w�dn�u�ν���q2"}0̅�Ȯ�Ŏ7)�a1�}`G���_�F���8��#��ʽ+�*��a���ZYHT�e3�T��&�y��������nr/��(���L>���?���dܪ&��{{xtp�?�D
v��z�r���X�f�q����u:���'h$���<=�1W�5�J���d�\��N��WA�Q��&T8  ���9��U����DOF
���o,a���0O�׋ՎkQ;7t�տ_"ܴU ��?d&a�,�vO�a��3��f>>��ܥ�K[��0�@A�ȟTAG�P)��ղ�Jn�}V/�޳��,���b��o�׽�a���G��y��"����0�����e��������j��H (a�5Y�k��k׎�kW���l���Z������.��l�og���1�GX<u&5���Ļ>E�f�8n���~���q;h'Ŀ�dHK������s��ֳ�a����[�\l�S�s ��^�B�)�8bW��هJ��d���`�x�pK��&����j}M$v�)t�^�\xZ�A�0?mk��|�x���Bv����{��d��SW<�Ί���j�wE]���?-���\5W�i�7堷,�S{}����OۭV���P]N�)z��Ke����Ef�>�/*�@6�b�}蕙��2~�X�E�-�T�2d���I9�;/i%pg��W6Z{���ɐ�tW�ۭ�[������l�vm�t�.g����c�-̺pJ�@�G	5.O���Nc&�<vs��G��	���S-!����d����D�$ꀈD �Ep�\�(�.�vf��9Ɣ�IC�j�ܦ�b�c*~<���S�K�ϳi��m3w���O�ryv �b�ē�F吼,���%�����M�����ߴ�Șk���:�G�y���0 �j�Q+��k%�F�e9Nk<b��_ìR���W����c�8���\4K������'费GHvA�c�{�z�0��-��EHЦZ#Qxc]��c��Oj{�/�ۃ�'g�ܝ�R�[9���lh^oP�
Ms�״ep!B R	�w��rW��p�E�Sd�._F5�9�u��L:'��ݪ719�j�%!��~���:�4�?�}�\y�0���!!��W��&+��\���e�8�:��·�cWKAuq��M������&q���k	�N���?���ڳ3Å���;˗WĒj�q��x�m����74t(�>:�d�������_q����s�S{��0R�/M���c����'����پP*�N�����S��'��Bx_վBZ��~�Ѱ "�h��%��5q����8�˃���	F���2��^�G+,���gyWg���yqov�7�u\� "v�.����3�.�Iύ^ �Ʉ�F��Tq�o���&���>��zH{R���~F���/l�������ȕ�Ґ"e}}��el��h�N� :;Tio,+���l������*�!�k��\�p�^��`�3�β���]�p�ޖ/����_��Ap��J7��D�?�_� d��LG�׉^B���]�Y0ՙC]1�p��m��j���7j@B��5eu!Y�n�+�o��z��A��X��Ύn��q'z��e����+���Υ4�����8G]�~��ڵ��޶9�� A�u>O��Xf�)�����Lb�T�+|KZ���]������]���A3t�������?�w���C���P`ah'q�q����曚�+H�DD�r���>,�륓���+.M�%ڲ���)Z�����	�DT���h��H�h�k/�5j .��������e�m]돓k
��k���K`�׽��݈ژ�?����X��pVst����M���8R�Cu1���?9MG���umi�z��=�Me�]OW��D���/������Cd����S��T�J�U�@/p�xg��ϒ�r�z�t�qp�0fY꺜�J�w�I;łj��2�,ɛ%A��ߚ�c�-���c su�P��Eu�6������}[���U���{̦+_��f_���w�v��F��hÄ��ُ��cX�I3s���&"s�w�~��Ï~���_/ٍ�g����#0��xw9���GIτ��zj9 �%����J9�Y�T|lf������%�7���HhxT�[/+j��I�:^/����E_s�'� ݘ����G(!���m�ҹ�����4�^���z���=���v�6[�b�?��/��������-�E �o��C���V�
���N�}��$˥E���e]�O���L����(d�y�^R�v.Y5�}څS�?4��m^g�Q��d��*�W?f�α�
�s",�����r9�T��n6P���M`�*���g9p�wDe��� �s�Q
�ץ�n`�g^�Y��|Dz^߷�t`��9�bፅ�4�p|-|7�)�?v���ݫ�k~G�f���'>���u��m˂"<c��s�O�����.߲}���y��v�X�I�ǚ��$"ʘ����h�\@�Y��;����_����U�3D����;�A�����KW�\� +o�[���PB����"�c�%cs](���-��� �v����1�KX�@�^q7O��
�%11d)�~�@�Ɏo�����s/�������y���6�E��_�6�J�P��?1q`9���cYbD��Q�>r"ɘ�0C�����i�!�-��;?90~x\�6�(=W�Tc�mceP�G�*����4�!���1E~��dVG��B�,bQFU�I4��@U�(�+JR�b���E.�KR� K@��(�@
&��jTDPF)�l�
���Kh�A@EAS�h|{�,QU$?~�2�ל��;����������O�}u~�?gE����@Yƥ�L*�E,QA(���F���������l��������h!c�?�Ó� ��'���~�+?iWM��s�Q@�w]���E�!�w\�T���?s\�ϛ%>L#��7�_�KV����`u_��X����M>��%�
�#��&Ql���%=��f��A���|��HM!�S��1�C�N#�t�1¦�7"�6�0���,�±�'�����V���ц��[�1��?6.���QD�%]v��/�R8î%Y��ZHCq<�}���~~��>߱���}^�}-�a�!w����@����O�;��<q��_�|������$�x�c��r�CW�����+�wF��ה�.��\���cJ�vF�9d��jME4:��Q�\��P�v\�9a�]���k�r0��Y��g��ڈc�o�g��{b�a��,M:je��j����j��d��&���ݑqW��\����?Ƚ�`ּ��j=9~ӭ���`�/�=t�̻?��g�3j��>흣���dl~ե���-+n&��`���S���n\;��$��1d�ח��p!��y��o�o������z��!U���.�����L/�u����~����@�z��p��#�D:�
z*Ռ�mT��N�����F�B�T�O!]3Qs��n�)lo����_��h�ũ��_�^��j�g���w��i�A��>�J��=���)�/N�(�ZɶR�_tSDE`�]9�������*�i8(dև<�S\8 宆�+��	C"A��H��ԧtԡ�/x��T5P�0Eb��Ɇ@��"�J�`������J��rd!�=�*���]��7���۶�ˬ���W��Q��O��	�y�?���ԫ�J��w�1­l���sQC��+����G0�</'�[���+��y��o7��Z���!������k� ����ֵqik%�V�TO�SL#�2�7qy
u��R!6��Y6V����_�0����ؑ�4�HI����>��=Y�|���,�a�!��&�/t�Gv����T���j�8#C'G���O����D�	����}�1^_}����%G��p(X>һo�̇����S�׼���k°\�.���o�얨
ó�U�PvL��9u2����%F���R�3<L�~�]��줒SD�ǉ[ъ{�s\W��h�.;{�����R�kWkWq~��|_/��|f�0cj��rO���y|����&���ڗk��C�j<�ۻ�s33��C*�N����'���轹|��%sPT� ��;�{�t���7��'=�^���|; �Y�{O˽$��c� ��!�B#!��k��0�$w��У_[��7���_���G�~3��?WiNT��s�$���4�;̺��I=�������ʶߑ��K�wӎ�s����n\�e�Z�����<�Κtw���=�?�f�ٝ��T/C0K� .��Q��J��@ NFݨ4a���3J�>�`�ҫ$�W��{Q~���e_v���oQpl�sQ���f8s�`��KQ��o�=ĸ�r-�u����"J��	�y�"A�}6[�LM�����t���5�LzU��"�"�̩B��(d^I��]�P�7z�V"������_��CD&~����\����M�B>�t> P�8:B(�]�*HLT�s\zN|���	�1�*H��3�Mάh�����b�1���=չ}ȋ�����C�X��0V�) C`J.�ymr"��y`?�9��p��xC��ע<�:�B����̏�=x�x� �"�P��Bd�.`SR�M�R���%0 )~0�" �`���$���*���P�$����c'�|*�D�,��HV�J�Q#Z@@��%��Adb��)���_~�7��NO0��)���UnI]�9�OV��P
R�Y��3ˮ�pwB����~��\ѯ�h�0�d���GVگ�X���]��:9����m^�V�����ش���༡�Ķ������k6+0��]��Ta����
'����8)��7�>ո����`�W��5��_�U������:��d&g4u#.��}b�[�/�_�r��1�Nz���ě��s���S�O��;�B;����h�}��v����zJ�ׅؒ] ,��7�}I�R�1��ϭ�dB���[_���w{�8q�ĸ��l3b֥+!fg�J�0�}�.fbOLӊ�a��û?E�m{?���_vk� @�`>�����p7��j��P+)���::	i�Cd2�!��f3o�pPE�"��,%���Fl����UX0�ES��j6��!��X�W���[2�����f`2\�ā�w�)�S���[ecE���h�T==2�����T?%ϥ�D�B�hd`!CT�\�=�3�]u���>��eؓn<�l����[��/�<�G��Ny'#O^�X¡���f|��X���$�����?���]���4K$�s����x�P�GJ,F��B��" �ɛ&<XO K-�SD�+]�T�ص�8�o`rY����9�)e����o�P��PD$ ����^H�,�! ����tG]�rq�G�~���;��''s�;-��0u�;f�UEBJ%%��hss���\_�{�B/��cLdL�/r�����=�]��/�rծ�MO�	�5_T2�*	c1��l�U��|�\f��D8 ݹVol_���.'R�-�+1�t�]�$����g�8|����~���������2���x�۸!�W�RG�g���).FA��d���?�o�~��eOG�}G�{?�xi�}�z,Z�P90$V@�� +@��l-�{j���aLn�ū��ק��� �J _��ve<,5,0g������ڭg\|�e��^����(��;)L@����B�A���"��* #��/�ry�g�rm��1$(�yO��L�b���g��1��V���?-4l��e�-�q� ��(@U�,�"�H*[�۫�8z:|�}<8i��b`���Ğ˫��u��:ov����T;�������e���Ȧ�Gj, �����Fl�!"wzU'Us]�C�|W��`e#�e���z���)���ֽ_��2	A�X ��]��uܶ^������,�i��u]}���8�	��.�k�������CF��o���I��-*q���?gBe�J�E�hH���=3?g�a0�&sWV�7�/F[(ak8S��8�ӆ��#a F"�+\޹P .���d~��QU������4��:�K��6���Jҹ���ߑYu�sؓcO��@D�X�m���돃�� l�(�PAއ""<M�ڭ]��O=�
���x;&δ��M*TUu�L=�e-��.H�F������׬�͎&9��F�`�JqHM黯i��0�srh��� 0dDC�����YX@ �A�Ze��]����� h���4�&Ӯ��	��1,���!��o�br4,��?��]�! A�����T�Բ���Y�����;BG�&U�c�K,���I���o2,(/�8ZU�_6Β��}uá*#łW���%!����p�X��t��h�6�w�fѐэ:	�Ī+��(��e��Ks}���h7�U��N�����cy���rōb�W,d|� ˫�$ �}�ϻ���t��΢�Ǟ@ȍ=?w:ő?b�Cy��L"Rp�'�zm��9���|�Y��J���BA]���[���B��5�`����"Y�h��w�fB��s�$�6w8X`	�`C�d�c��,�M9lc԰�������*RBP��������maM���#���F1�D��0H��B�� �X�mJ"=)��a�7�\��"?����3l�w�ki�����-��������#���ﮑ��}_��9��G섵w~� }�y�c�4C�����������w{}0�G�#Id�{b?��ZGz�>�>�?��N�A�G��j�nᏍ�� >�����y.C��[�ΣU��!~�[���ͽ����׈W��o>>B�|�(���9ә �S��Ԕ�x�a`k=Z�2q�@c����M����p��@��	�?TT��p�3�%�����5�^���9���;�.����l��Ng�N�~^�ZK�<�&��}k�}�	�xG�3&�L��=�B\�����LuKӒ|]��jl9���hS)cD�*��XX��dI>v��h�*�
��&Nmُ٠fX,R��)�\�����;{ꙩ�}4Cf����okc��Xb_c�����6sp�g��{���ѥ~�c��m�q�\�ƇA��G=�_C��S�! ��;�x<yq��|H�|����u��p��jF�P�D�PT��J���Sy��k d�{�s�ڻ9��|�'kSK֨�_����@����Y��|v|�KA�`E?3l����m�J��3�Mn�>��d車��q1봙K�[f�!�t�,��YL=&k�B���y�F�M�C,�z�ꚳ��ik�@��/��V�a���=@��B�O*kz���3�^�,��wXfk�����o�Sa��<��=����y4�z�_�흮C�/��bg��`�����ԧ����T��iiz�~��uJd�&�=j��v���j`>��c�"�Wzvb>��y3x�Oo��|�J�:������,7K���l���:>��pa��K���N����[�"k��tC�@G����(�=�F�j:�����_�`���m��Vf���RG0%:��3|���y�T=2W9�|k:|�8�R��ԁ�g���٪<����r�&u���5��l�_
��ck�t�\KP�:5䬧Y�����GW�?q��p���N�A `[:�}���+X������:(*)���P���ZP� �-		�@�&����Re״._v���a�FL}�j���S�캼Qua3��&Ad!��lH�Im��%jQJ��)B�a`@��������+�?���~��G�"*!È�g�	D��(TR@IADBDF@RET�$dED@UdQFARDd-Ѧ$xUa9���XHȩ�����}{(�!�a����+@�$�B@$@UT�"q�[k�r�U@x1(����A�� ��ٯ[��4h����XD�@B 
�! ������q8��T5�!�cFn�'<U�����^]s>|�}?N��zTMu�w $����oH�>/�H�x.��T�S���0ԇ��ϙaA����[���v�Iް(
>��T�T KV��"��0bA� e��q��@� L�\�$J�&�A�D�O�"�	��4A�{�=�����?�����6��P׈k,1bE�,��!�G�� �m���ǰ" A��!e��A��шzG�����{x�W�P:&%@w���a? ���"�� ���M݆�E���t@|?u@=4w� MS����3�ð���a�A)$�@$&x.�G����X{��m��H8��L�����ͩ����R��(��дՎ�]uB7]t+ݣ������FO<H�֙�b"d3Y͛1}]��)�.�2#�l�f�����JA��Ĵ��-�Z3�NO�2�t���A�Hf��x?7�ƻ�����>�&x�g#E �b
4�� 3��n��C68�c�<h���͛6b���
�C&L�����q�]Q�Jf"�G4F�F|ٱ{8�2a��1p�a�����0��#�a����r�Lq����L0�$L�lq��bb��h���wZ������Ns)J��e9�e�c�-`$�@���U
��!�����:�?Y�P�j]t��p����҈�P�1�X��y�!&�������qf�$���u�	 Ess�3f�ٳ�I9��eYe\8���,�W�����{]^M�n؋�0L��ۡ��
/u���`0m��� 7�?_ i�W��޿Z�Y�Knʓ��7R,���,�õ��BKL�T��4���^9�C�r�8v����� ������,�%�Z4V�����f f͛6\���c�$S\/�����f�����U>�C��m]ju�<��1�X�X�����(�j񙌹L�/az��t8a�K��
@c��7�F_�=\�ƌq(�����_6���Bꁢ�M���CA HA&�,�\6��k����P�#��#&�iH&�q0bҠz�3v���s~c��듑��cd�̓�u0�vĆ.ڔ�,�9L�0je�Y�L�Ø�ü��iV��+D�D41k��v�K0�l�b fflb�7vG6<��~_�����cU���ξ��G�?q����/�۶��n����I��˖��P�ٳ�9��xJֆ� u�	�y/ry!����@!�b'��A w����K,��@oA2A"qAd����|��׻m�s~Əy��o�2��=���c�~��@������kPF"b�h����|����`��C§�Q?*u���'�Oe>d�)�Oi?�����'�O�?������O��=��I���'̘�x��@�������ĲA_!�=����O���$�S�M�m�n�t�������?B}����'���<D��M:T��}���y=�?'����Q�#��������b����xffd$�W�R1Jb��N)8����^����������O��n6�}�~&���Ēf{s����I�YF�#`���0���������r�;++%� `���ɔ��@��Ё���9��9��9��K���΃��6��3�2�իV�Z�������X0`�������^���=�>;�PQ_�JH�H��^�z��� �.\��ݻv�˷~��s@����pg���~Dp<yb{r*�*�=5� ���򠠠�ſ׃7u]��^/���pv�������jjjjjjj�*�P�B�U
�T*�P�B�]��K�����������!���ǈt�p�eG�ٔ z��������aZ����V�х�\.�!��G��
���p8�q���:�a.
L(
p{���]��AsF]����� �f�!aQ��!�1��.F�g�٫��x�����|���;�y��?�����G������h] #ނ:c�R'��^�������)Ԧ�J�pb~����55555550_���Ӡ 鏔�����t�])Κ����w�������>׵3��+���t}Jʀc�9yt������)�11.%����P���F�$	����{���lW`�x� ��c���h���jEv�}��o��������o�����}��/����uu�/Ϛ���a��}�U��1}�B��`'g;9��5�d�/
]��Uv:���[�� 
�4e�]b��o)�R��k��~�R�_�_�&��Xu�������V��^*����*��XeY[[[[[[[[[[[ZҶ���"���K�Y؋݊�iB�dCx���UU.�:� ��[�`�x4�^��^¢��c�U�*�%�n,V�⨾+Z��&��#s���w;��U���R�������(�bqi�N12�L�Z�t�������U �W�*d6�G---+-'&$���ddd䤰@��Zq�9�ϛ6l�sgp��$���������Z�v@s�0`���+8p0>�!�H@ u "@D82y<�O'�l2)�F4��)�~jo���fff&��**"�����������j����{A���S�y'��\�S��L��rHrIɜ�P;0Q��2�"2�{Ǳ�O0�i��Ye8 /��d]|Ʋ��fD H�U��P�B�  ( ��? ��t�Z:�A�kՀdrd2b`�A�=��-�FW�1���9oj{Zͥ�V�ׯ�i�O����=�}�xx<�GC��9�u�ñ��J	�L�2C�T<�TTTTTh�z=��G����z=�G����z8"�.�t��]"�H�E�.��������������������������7�?���?��gغ2і��e�-i
MMMMMeUUUP�dB�Ȉ������W�}��}���N8�8���'Rk6�M:� 5� $� ��o�jjj^jf�'�﻽�Wc[ZA@8��z���e��������N&�M0�yL���~�R����3��g�(������Z$��|	��YP\S_\��kMd	�E#���Z E����e�=�ǭn�8�m�R�*��Ɲ��r��~�>�\{[�T�}��{�zݨ�xy	�|��M&� {D�OA�,5t��!��$����i\q������-�]�,I��,�縊��
�WQX:)q�Q���2ry''VVdKĤL���>9��s���=��g����{=��{����w^�	0 �`�t�;nz.2��@��m��D1��0H�@��;Ȩf����|��?/�c�ZC�ղʊ�@�R	Q6"jp����~_i�9�C�AҚ ��YLS���O��Ĺx�* , ~���6�P�}#�q�g��Z?��)�flc&�3$�@���-�ե���	G��6�L��VQ�, ��I�p�**
8)CL ��m`� Ȅ" oRN%����#h����H��.�"� Uxq$!� )�@3�st]E�t]E�x�ã�O!���@"�T ;$���)m?�6��ՙ�	|jz|��c%	5drfB7�	\�!���H��ۙ���x��C)1���M�����X)�h�
��&PL�u�����'�``ɰ$�D`�C���Xq1Z� ��g� 	"e� BaQN� D���	B ��m���nUs��闭��Q!	����/���E�5��-1�\���\
�����A�`�4���PR�+�%ԃ���Q�j�w�� ����r}֗m{�͝UsHbo{��G��Um��a��U5�6���?:5d��iׄ��`����}T��Y�n�y��`B�u1O���}_��c��>,����?�g����|��[��}� D@Ȉ	� �@�������?Ӽ����3�S�~w"�[��L{��yڋ��M�.d���t�����'uڞ����_��zz i�B���oD�J�����S�8�S �C�wv���H�x(�A�t��.ۡ���kZ)J�@�%5mDy9�L��ǖm�4��fه(vVO�����ivt�n��
RJ"Q���K���T�V������hq��i��^-�/���HBq�a�+�����e�]҉�\8s-i���z�^�F�u��J��kT�j�kz�(6�橂�S(�R����͉�ް��V��j��خ%BX�^�)D�QR���/(I��-�f���˵�8A�aS�,�!(RD���ӽL8I��2N�SD��]���̶ۼ�r��i�xv��\��ը���Ì�6��7��Bu��8��:֜�ckAE����]�+�h�5���������b�6�em��1�Q��h��2�Yn��SKi�f�f�j��Q�4���pۅ16"���Y��	sNA��Ѫk5�e1ۭQukj;B��w:f�oa�N[ےn�[�B�0 �qJ�.cVSTK�R���!	Q�.��LL�tU�f�Z"-K��5�R�a�:պ*c�j�wscLfjeA��F�e�Xp�ќ����F�(jq�eK�Z����B��֕ۻ�]W�K�x��	�r�-�m-��LsP�m�\����˻8�ik5�
e�ZM5�m�\^2�5v������T+�\R�T˒�Z�tj�
�� "�[�w;���$� �� 6�b(�H���# �D�� �7V���oÛ�Ry�i:1i'N-=>��hxP� �������ާ���{i̥�=���N�����OY=d����o��'"�����L�r��'���TC� ��# E	�����<���Ze�<>.�֜��Ɗp���٫����:77u��P��)f*�xַ���jT��k0�e���n;�a��.�Ùr�p��ȨL@J]���49*]w5�q���v��5m�1S�n:0�T]&+5e7%�V�]�.�������x���2�ݱ^�QA/����MU��a�k0TG�B��h��L�.qnj�1��kW&*gK��4�˲�em'����jU+�M�یL�ư��-�G4<at�Y�*�5�b2�6�p�Zķ���83Y�t�4��ven�sJ�O6�LN0���3�#��Į��w�R��U�f��W{�f�b�ۙWv���jQ�im�wCN�n��6���Z��sF����\qZ�7*��)m��k͙�:�R�UD�&�8����ޱpPkn3�Z�W�U2�5Q�P��Lh�����`�<P��j����s3�S+�tYUY�Qu�Jӆ�fԶ�.�oZ��]���*����\km���1Eƺmn	���Tq�6qnp�`�\��wY5R�w1x�L�,��f�f��koց�%���+��n����0S��YV��im�n`�X��]4�eʙC*;�b.Z*�qf��c�Tި&4���h�ER���\r۬����q�1J��E��`i1���h��kG.dhҵ
3�%�N�2���-�ֵ�8�]1T��raiU]�*7[��A��d���tԙ��j!*��9���1w�\pv)��cX�ue1����콄�T�ΥlWee��s��� �ɮmk�\�,�_J��]G.��n�<ݕ��o�rݻ�ѓO�����k*T8�S|��e�Zf�ց�6�Kij�i��k���w��s[�<h����:�9 ��8A���+�9>fO}C(�6������R�@U�K���Oc�=�[��h������k��k[;�Yfu�m_��o��؇��Q�<��Z�W
��@�0Q梿3�s4}� bxӛ��܃~p�ࢪ�Q�@j"TU�*5cc��߉�o��Y�����D1�6OѰ2��ޮ��o�ߤ���X�ʾ0w�>��g|P Dp���(r�U;^~���U}���.|iB��Z"���Nv"#���|�q��ϛ�>�����I$���[M��
�*����n��)d�\�@�̈Θ �c�f�(+���27!�)�@=�G��/_�zH·�:����R#" �0@��<�J�D�5ƞ��+xE�킕H�2��9�\�.�
�s���U=���9�̳�b��ӭ�e[���Ph.��<	�؀J�E�����og:H��X�Yh"x-��`�	�4&H� �X\��n&&�T
?(�l"vR�$4y��#[�:q�m�~
����q���"�v;.����|��>o���|��D%��?7�S�'� �����Ƞ�R��[�tݚ Y�!R�Q��A@be1R8�/H���R�p��5cV����[�A<d����!��S$�D }x��DS���сx�c��ƫ Ȁ��PD@s!�gn�q��*����(���R{������)h��D�c���4th����@ŏ=�}(��G[c��m����o���z{��v�+ȐwP��d��>���5?��j�O��u�3��S��ޫ��GgJ�.�.���i�RݥbU�vk��:���Bމխ��{���q˺ϰf���1+�
ߴ�;J���孍Wc�+�2m!>�S�$�ֲ�-T���jXuk��3Ňk.�[�o��R��Co���`U��#�
��ѽfL�5�v]f�qp�[&�i+on^�܃��-͟/��qV�Z��ͳf��8�܇&�M{F���8,Z���Ƿ��v��_po�L+�1�v���
�'bYl �e�P���O��=�����}�&~7E��j���'���H�n�=���$b���0�B�P�����&�� ćи�s��_CP��Nv��vO�<���y���8�pwhi�t�$E=���]o����·���>�H��Ǿ�b(��cd$DGb"���G��~�����_��}�u�Y]��ځ�{��k|�0\�HDB<LU?��}��{�����/��������l y������G(�j
�A�41;~}���|?�z�s�gt�5n�b@�����9R \��غc�ֹ�ޒC���M^������
��s���$VO�eѮܙ�̝Ŷ%�����3���u�};7/x�c�p��Ya�.VuV���S����޵���аbӟ%d�/���+߶��`K�3u�p������%}�o�Y�},�՗*����n�W��V&F+�Z�h�I���v��*@����(���n[�����O�o��g�?�F^hXߦ�9'5�+�-O$6k��l��ar�*SA�k�@��eɹ�ŉsw&���������Z$*u��m׶j�����z�Lr�;���z��n�l�l�k9T�rf�2}~�Y���l���4E������~���V���5E&+�7"���y��6�w��*ִ��|�Z+d���<��y���;��q��-�K��ܗ<�j[�57�K�32�3�As��RaG@ @"��J� �WP����ex�  $� ����_��{ݭ�wF�޿�n=�3� ���a$)d�" �6�p�1o�������P�a�����^����~��<Ns�}�:s�y،�C$3��ߍ�}��)ek���U�>��d�A�'���<�_�c��F�������w�� ���?���T�^���y��_*(l͙���E80DC�~e(v�;D�P�
���A�]��7�?���gԷ��x���_�xܖ;��ᬱ�ܖ^.�9��DH0sh fF���A
�f`�ȉZk_A��.����l� �XQ��4'�љ�קcd����c�i������(�*yP�N�uS���:]���C��鴺hXB(�16�� �><��� �����o�7��� ��Z@^��>(�����g�̟*�0���1����O�>���j�Y!$W�}���G7���ѵ���*�Z�˭tڃO۞�?���D;��:������������)9�ϵ��q%�|�5<��r���>��}.��Y�)}�3�a\�����9Gߏ����4�O���t|�@!��&O;�)B
�.G�
b'N�O9�{���j�����`]:=>=1r~��x=�{��<��÷��O$��y<�O'����MMY���U��<+,!!
#C y����
��W��"�b�.y |�!����B�����iz��v�۶�ضrJ�}�M �c$F`|AkA�~O��v?N� �$E�mZ�Z�h-Z�[��'�yQ���t%NF\/�ϨMh�b�J�w�^~��G��rH�n���C�}%'�<?�p��ھ�i�K��J}�3�9���,<��8��ax��y�|J��o�Îs�y�����p�S
��JF'��jz���\�K�E���<�+����x"6q�� ��� ������_ګ�Ԍ^�ۿ��(A]��Owy�S�+�Z[�Iٌ`�����T*/S��Nt[�t��g|��������^�
��a|7c�1��cm�ڬ&�^HH���ޞX�o����8wg�����G_��O:���q� 7��3"׍���-j�v]T�q��y~�v��/AV:>Aw)q�"(|n��dI�6!�";Sgk�4����5zM�C�8�|���/�8�Y�C6w����]0B�X�������EH����jY C>�o������Fdf-�=�|�AW�F� �0D�&�m4�v!�X����a-p0*�n�0۶�޸fv�D�dc�I�� ݈���g\�;[[Yv����ǟ����,�US�9�������F_�hM2�(
Pԋ������N�ζ}��vg�z�F�]��ő�zuK������_6��������l����$]L�r# :��P\�U���	EW��2���d��Q(�����咏��'Zu'�{S��ⱘ»����7�_�n}�����>������L��9K��a# ��
��!QrQ Ȍ.)2D�C�������}����x0>�W��}�~��i��}]��������������2Ā�j�
M2��	  �� ��@P�KA���s?��M��i���!�Y.@�G���z����l���=�a�<?%"���p�h�"�<�������D�+C�T��̍܌��GO��,4X��րdaBA�Y��!��ah\a�����E�)�t3BҴ�j� ;}�Pfe ���i2���oe#���oe7ǩ��u7�����醧S�������ji"�Hn���yT���<�� 
�8�H̔	��ޭK1<(�^ߨ��
#1�:5��ц`� d �0(��h���������6#`a`l\�.{�������#����ި|s68�m��3�?��?'����19s�R(P�s\3[WWWwwo��TV��ֈH����o� �c�������A���@�P��j&�{�����������κ�ֺ���",DU%���شE��N-8��S�N8�Kt�X����J$��7�h�`k�)L�ʖrrlV��!��`�(1��nnE"�ʞ�@�!#"$aiȈL!������v�Ev�qd�d�b�*�ر���y��9�sy��9��o7,B����"�x"�8�ē���0��|1;�YOYYYX�T�.�/:vޒߝ��C=�P<�C��@x>7����@�B���Dexx!�c4&�'G}�ڃ*��|� ���@Ɵw+��z˾�?�P
�QQ��C�R�\��{%�`���;�9��̭8+��}����F2r�b�oF
?/�Ӣ;��D(�$)�#z�a�8�Jf�9�=%8c���k�{�ξ�Е/��!o`�!$�?�Jm4�+[Db����BN���m��DD��Ϟ@# `"l �d�tfXo
�X��p�����o�jݞӗΛWO@�]Ҹ��c���6 ����"�jD����_?�yѧ7�n8
Z��n`1 0X �k?\�33�U�.g�{6lٳI����ٮ,3f�VN#4�iBJ�ǛC�f�x4G��X;5uy�c�9��=?�䅍i|d�(Ȋ�l��_]m}}}}}}|����u��W5�������^Ν~���� kL��^� �Oe�q��ʀB0v�\���Hdrr�uW��n��q��l�G.I�9'�rMsXA�J-�a�k
)�ލ$������ϑ�@��� ��×�I3F�u��� 8.�wCV^���1���&�"a�}vW�ZA����q7I8���[�/��F�Z�Z�:�9�DjBg��˗Q���!Hid���
���O?T��:{�I��$�\��&㘩j� �Z�7���}���Oll=�^LX�HŊ=�����d�z�A���"�>�m��3��t{�t�iω��̈́�y�r�su����.@!]PS@X�s��BPiA4K�\��Dam��9j֡{/S����l��:M�#WFgҧI���,�N-85бv���`��߬i1&C�<�O��e�s���������B'aԇ3Lկ��3d� ��I0��:"J\�v�HA���nw�x��̦&٤�I���o���K9�����8[� �P!������w{{{����޾G3�ѝa�q�Ws�}FV���/sԖ�ip���_�é`rh�u�f�CP�sF�*�M2
i�Ʃ�$��	/Q�F��A�f@NHA x��́4�M3�	���И>
%
�ddD���A�'��e,A ,|h�@�C�!==�(���������$����0�� �c�xk�d��+��P͑f͑f��l�͛6G����|��_�5  ����G>�=g�8p������-A�:=ԑ◄�����=J<`@G��O�Vl�6l�6l٦�f�&"�����"#`~���|�g�p�Z�D���^3jTzY$���UU
���E4�P|@@�`Q���V	4��?�R�sͩ�-��?F��Rw/T	@ςIׅ�ׅ�׭��^�"�zK&��X�A�x¨�i�	�	/Դ/�]�|ҒH�N�k�� �T~�nx�8�X��lbŋ�pp��4 ��u�m�ޛA�X����нB�c@B�#0=8� �!��~�����/������Xch�a7@J
�	 kѡ��X��ie�V1ƽ��飠l�_GΚ�r�5g�g�4���'��͟8ϟ5��>���k! �4�_��Ӊ�`ы/���xt�Gû�i�1X+�"%�I'G��q�2G�H� � +�|�IN|��q�>l��|� ��|h�2�G�V���p��*<]�<�>h�z	�9N����4�	p��M`,�tY��|.?A=%~��RN����HV.�o���h�ӷ��~�3-��QQ	I��fzvrxI��0��&R. 5$	�� J$1�I��KiJR�[F���_->�^�����1,�:�7� u	RĞEm��̋=�b*�S����]���f 0v�+��b�C[m���Tk'*���D�d���U[j���XD��t�!ŋ`Cw�$SA5A�,����ȱa*����V,YR*����
�� ��!��� 8N/�~E�}�<��I�s�URUUA�4t �N�H��u�1������1	� QvE�q��R17wuwwwL|�W��.RO�!C��www�M��� mID�4�h!m�`�o. !0�D#\Š�%�X0DZH+�pbs���\3�g�Xzئ8�C�Os���ls�vI�E��KcJ���'0t��l�L9�)��K<h���3�������K;:�z=
��&� �=e�[��3pp��CS��p�5`�^aJ7t��+�ժ��y���Ǧ�-wP�:�%�eb�?��vAv�d#���W�~ف�5G#�ߦ*�A�"rh����sQr�W=�W6�M ��!b�>������oAKzxp� :Bg)�qw[Cj�b��d�%%\ �� ?N�mez��|6�������L�i�
���/�0����P<30ݿ��}F��C0W$!�'U������S��
��������������ԐT9��G���Nr9G#��Mr���P"�>����!b(���Wn��猃�1�D@��fB誧�UT�˲Dň�E�-	�$�,�������YD���81�_����}4xL;��	UT��-&��oii�Q��^�|�x�C� s"��������n7��'0[=>s���w7����ӝ��O��� '1�0w�0E�H������щ;�=էm���f���"�$Am� e��"o%A@o8�^�"v&���ǚ���4:%^�!ܥe�6w7=/��=5S�!5C2u�@�ǯ�B,ºJ�VR�,�*dC� V~�xp�tf��8Tn��0(�8+gd��.���)�	��Oxt�dn+6(�6ut�5rbJ�$�ӧ^����^��B��5���5�|p<uuh�@���=���F�� e�S�Z˲�VDA>��Ӥ�Ś�,��9����Ϝϟ?FdB	 .A�l��e�ԀA�F ����nx����_�C��z�ۆ�;dY���[�o��hkh��NfL�V��?�4᫩X����f�:�,2!�~���5���(�HD�3)�l^��%�����P
�nDhHCs��:��h^�����7��ff0TQd��ՙ !M��SY�(c��g"+"�8sN�I�6�����E&�/��QȅN�=�
"��m�|���	�nh,�"l����ΆL6�l����p@�u�]��Н���Ȱ�j����|��/sjd775��ss�v���D��㨁Q���mP8������Ň�¡��
{1{\�'|��(��ctՇ����9~N��� 3��� �>�p�Vڜ��U'�öw ��£����[�ʦtѰjeI1���+J��篕.��RE� ��7�:�N����{>�t�7���^^g�����Y�1���vo������Gw��D�"��	Oc������:6�
�@:P<�=�U��*��o[������v(f��6urn��>�J'�J�(�O����N�\(s�z�~	o��E���O��x���q�p�~~�Ǎ$�`�ݑ���T�8+P�瀪���V!΄]��0��?"���|X�DY��!���G
��:�O<�'�$�C���>����o[����*��!#)���r�3�|݅��Õ�W9U��9�%�H�m� lO��������B���f��u/#����Ǯ$�__�\��d%J�*�XR��<>��?�x*� p����QUQUVBt#$;�����o��9H1"���͛�7&�;��C
f�%���0"*UE���Ab�����EF���"�tVɳ��m�֡�7����}Zey�(�8[������c��N.O����-����=~�k�Ίh� �98 ��H�*`�Eg����3){T��y�e**���,X�EQb���(��)EQE�AAb��Q�!B�����x�=8���3P�U
H�=P@���8t]}���I �ߕ'_x��/��ֆJ͛x�7��A�r�a $`���mcJ���̧j۠�����FTB�L�Ml�ѬkqqI�(y�I�A ���g��WQ�^����y):fo�<ƫ>���+��Nv��Gk|	������=\2(
(�:f�j�	�r ��{�����6����<��=Fp0�4f���m]sR�l����BF��$:��§J@0�
LI�M�n���m��\s���]h�Q'�O�{}��_���>����r���9�������ˉx��`�*j�U��Ut�ʪR�L�����ʷ���D�$��c���u��/�c�e���� h��y�\��Х��//Y��֪�p�ԍG�i��f����۹)����HYK����щO�~���&��R��dq<2�\�^c�BCos�Ye�� ��Ŋ��e� ����H���K�ڷy�\��%��2h12sP$�	��1��t$��属S7u���}��z�~�����:**	YZ
*!�y��U�Օ���%��s{��?ɩ)�B
d�Z�"EWpEƄ�,�s�LG��L������j�R|W�h���a�T�Rͳ�������������=ى�����(���F0����|#�X�����İ����4K��L�E1���w5Z���[[H��V���|��Fs�K��������ώ.�xxxh��uW��[1�z�0��X�&M@{���Z �@_�\�A=�uTν)���!�t�.A��~����L��	�D�d|������������6$f�������~�y�ﺛu\	k]�ËX�B�e���+}�8�@ R� 
`�	�	�������5߰�?^\����K�1Ď�{��ݻ�g��Ǭk2�m�NA��F�qb��̐E�w�A		�V�5@{��Ӵ�,�@5��Y�'��G�o!�_ p�2c�����m��d�s�g�
��� C�ŝ a,�*��%(��7cT*N.���@	VL�u~x�m��m��m�m��m�71�a�a�a�a~�b��I�a(+`ŀ��p"h�P_�/՗�w��y�hw=By�zIš3E��98����!x&G�t̂ �ĉ���)����|�F�� ѱNx���D-�:""c V07�H֨�wwv�!��d�R�?k�����wW�����8��9�3Y���`)�B�"��$���%�/���ks�?�f//,������PX��0
�6�k��|sX�:}}|���z!�3~d:��`��F���6��aL���6�M��˹�e������y�D�m! �.��ˆ'Ə�3�C��X�bA�b������u���t�"�<m`)����";��O_	9m���>N/��0?S#��`#`=����Ȋ5]�x�ð��81 ]�H!Rm�����NIh�8&Yր�������5�:�� (�~Aڂ ��@X������04����'S3 #LM�tC�w�����y���C���{������q=�o�;����I<���)@I��̀D�X%�P���KMQp�?g���{=��g����|>�����y<��U����~@D}�B�d~�Ǔ���y�E��D�ȣl�P(�YR��A����EAT��\�����X}+�\.8��dMb�!]}0�2�����3~����������������K�z�}�Ǘ쨇y�s8SS�ȡ��vGG`�y��	��N��o��: �#k=lR�x�ޠ�̨�>��]T"O�A�X'$I�V���X>a�@޳c�n�z�4N0fb��"�OM	��)mZ7L�_�P����HȹFD@�}{8Sic�-�.��af��b�ac	�����~��o�y=֙�|��и[d�B�����A(G�>�G��]�p]�����d��^8?զJ��~������\�OS�:� �,a����pREP2��]�`Żv��l[�d����*BLD|�W��J�I�͈�������O'��߽r 4�����570��3A�A���2C!"A�z����i��N������ X֢=Ï}��g�8�F@����/��ϝ,�&�i����N�?HI����Dju! XT S���_M4��0]�䟫�kcW��O�--�%�rQ���F`���$:�����GZ���(�P�"6�	��`pl[o߉�Ѹ�2`�F���:n,ƛ�/ݼ��)O��@������[�Ʒ?�q����2��74v�Z�lzܯ���ÉD�"�P�@wtoI�xI���Ŧ� O��8˰p�5��r9��|�I�ϰ��(�1b���)���#�b�V�Yr �\�W�v��G�P�Ȁ��2M���)d�.'�x	c�������é˜�,!��q!�qUѩ��oq8�����<]��"���<�3�v�4rl��QEQEQEQEQE	OqE6�4A>�(�Q��m�ɶ�m�8m��jh^9��G�;]r��j�Ĥ���0��+$��H�&�q�G��w���unT�mD�UT+ ���ءT@A��Q2�ĺ�ZZZZ/ciMiih� ��7h(����$�<��|l���)UU��	��<�P��C�������he}́�zc²W-�잓���9�
��=�v��k�m՝���|����`%���wx?}7��-9�-��!b/��X�?�r���.ΔBN��9 ����U@��h���}*�wԳ��)5�L��dŀ��0���9l5r���aȀL y�����ַ����>�Խ����������
V�)�g��|�`v��~��0�n�p�V�P���ķ�p�x�d3xv,���������28ti�7���g�m�~���X3�tA`�a7'�z?��w��x�)�o���t�lR�dn��7�}�.�t���m���p&���������ԸX��|:�s�	ng���j�	�z^6�jn�f�sQ�mg�~��ZQ��^fEO������(;m#�s����:S��9�%��4ձQ��}=G��.JJ��_|�����S,�Qʴ:�p�i0��q �]	K��P�� ��2x$r2\�������Hx�(�I(ly��\�F�؁m}m]�^f�9)dt�zNR�g`I���Nؐ#�����L��������R�:����6Z�a�-"��铍
�8�� ����'[߼������˙ξ׺�z41C���������'���wW��r�um��3�Sf7"���s��ؚ
�.Hj}���a���lp�N)�Dkj�������i��."���5/x�|�K��j�U���9�rַS�B/�V�)��ԡN�ʺ����/���s��n|����0C��ƕ]��r٣UCDr[��=�w��H��o��w��W��}'6�p�q�!�������.��������}��	�E�z�!+~�t,L$ Z)ғ�-�kR���ޝ�F���0u����>��Ωhzn�u�]m�``F3�����Q��YC� f,b\�魵�ߦ�?�r�`���m�0� �R�)���$��Ka���Yt��]	A,��;�?��8ބ�� 2fdyLM���-6s�@��*���t���G������ �\e$� ��Zy{�
	"��	&Xj����@��e�iy�U֍sA{ɳf�}�2:G	��m W�tƭH �* �0��"���a5���ʝ���Cr P'�]9��Y�H����S�Ĥ���2�Wʪg��'�7x�8���=$a��?�<���{v9@"fcJ��$BG���~�e��#�3�Z�W=NQ���8�5j`~�D�>z�rGa�@!� �(`Ŝ$�m������y�{g9�*F�6k�{�#�_C3Y��\�lM0�ݩ�F���g]�`������i-N�GW�X��Ad1�`�pu����_5c���ه�� �ח;v��MU���@�:z󡪛%��ꉑ鲉mIĚ+�n�~��op�W�����(4XaY�KD>H��9$Z@�BB��:!C):�� �`�L��#���M4�M3,��H@m&D�&bQ4h�b �0�@��֑�$�I${�6�%��R�2��������S�̀����Ye��!)��`D���!%D 2�����+��,�� �ڕ�� #�uȄ�&\�e�v�i��dU�g�S��ĢU� �٘ `��998����ѡ:���>�D�-&��.Y+�_��KW�Bqaz��5|��u��WѪuMYR��-��SH�쾎v�˻d,��ѣS�v�����;~�E1����i�ݮ���<p���7�]ߵ>��<|�O����lya1�)�Q؇���*�����!3]u �^u����&O��vlb�xQ��Y,ې�ƿ�Ưk��xZǸ4h�r�� f��je˗�)`��$!������^����ӣsg��m&8ٳ^��Þs���cq�>�6׽��u3�.6AwYes����YـZ	�5~|�����s\�D�3ʘ �uއM�=�l��y?ZY���RuI�O��$ڧD�d�ӍNi1�LzcҢ#����3"0�e�@�  ���q`}���6�C��0��8�� )��*��F�����>��{O��i����3���%*�9sMx4���h��H��#�X �`���3�($46��x�������j���dD�N��Å�D�eL�᩟�
�2A��ߓ�����:N��������u���*.C�>߯:�a9���ާ\y
L����Ԗ#@���A�Yדf�Jٲ���h�f4j��$�{��f���Ri�VKt�4��i�˜�����U���ޓ��5�)S:J@uFBCN�A[Md����2
�_��{�a�]�e�C��Gv���[@!$����<ݻX���J L�r�ɒe��7-l6%&���"Z�Ad�.DȞ�ɲ220�,LsUI-|�FE-�V��#�h�k��Kd��%��庣��5K�6��ݻL(���h�[F�h4&�c�b7�Y65!�*�=��܁˪uL�I40��a*pp}�M�g�g_M��ȓE%D�Aic��h/�_�`����tr��x(�=�#������ޙ&\�Յ�z�"��DERK�sI���.ƵB�JP
�	y4W�g�0������d4h�����T�
th� iEa p�kE�{U&%%�5��`&	�@)U��Y������$ ��b��%n��C�ّf�Z���dD�L�.y`.AD�c�?-�O�Ǎ���=Q�+���W>�m����.ԥnR�l���X���y섹m�%`bbE�
I�*���	j%D�Y�Q���H  -T�P	@�EQ��* �$AE���h*T� p����E��QP*+h6��E�$��1�b11��LAb�)h �A[Z�-R���H0Aed1$�0���T��`J�Y�*cb-��t�"�+V�& ��hE6͸ʅ@Qg	7��]���S�un�����5]Z�qp�`n%��eu(�t�����]]m�0�6��Bb��sV�2�ۗ5+�M�a��e���;�"�̼%����1�Kn�f��U0ʹ֪\-ތ֝7Z�%�wn�z�Y�Ӊ���¼5t�k8��R��W+�T�+8e5xx]]
kNM�u�b�(�4���ox�Y��n��Wn(�7M.�♭Ax�յR��u��nfo36\�6�6�&f�2�FV-K(���M�⹚�[1.C�L֓8�M-�k�5G��x���`��c-�]�����j5�N3Y�q�.��vቋ��el��wF��8��0��IA+jk#lSf�qٳYw�"�j�V�0Z�hgN��xL�v�Ub���4��\̛e!�K�5���Ʀ�.e]j�k�U�Z���f�1-myph���3
�\�ͣi��oZ�4q�f��j��Ә���[V[U6���mZ�lvZ�ۗN���x�36j��%���m��ִ�)c�����Lxʊ��KkjȦ�Óf��ݣP�M5Ƙo7L�!�M*�A�<&/J`@�A�Q^���ծ���mr�e�ը��
����f��6T��9�ECN��Ʋm�i�i��uhu�XR)�6�)*ұ�mUE��5��P�R�KZ�F��3"0B3�O�sn.g���Š���#��=��:�_�������QD�4T�_ø��[�|kR��*��mV(Ѳ�j��UT`�~��"�JE ��E�QX�UA�-���b�k"̴�}�`"Z�/����=O����{ϧ�������o���l�S�:rJ���\��sQ�⮾��3˻��q��É��:�wEz�DF���̱�觱>{��_S��;f�8��;�	�#����x(3;	=���~"���?����!d�|�����K�^�0\�����=�f���0dt�`����'���;EJ;{GQ&D>|�k����[ Q�y�(3$e䥮��F]s�O�ɑ�����ϑ�)ND6_���#z����r`Y�����$���-���Ŗ{[�{}o�W}�r��������S�\��L>F�e�?����� =$ˊrR
�Z ��6�ڠ�������.Y�A�|S¡�U1��]9��-��=�P�\�Ie-n���-^���{~�k* �t�S�����z�EE�-v#c�x�����|�	���DΞ�|S����>HߦI@����L%��g�Wu�z&�%�O'��pn��>Oگ�W�'㞡�z���s菜W��O����r���]+lB��gNw߬��� �=�r�����>�q�Gܮ�\�8��M�
���h�?�_��_Ay{���<�����f2�)?W�B���B��*dC&e�R|[އ����\�~j*��;� !��Qq7��K��=o�����yz��O����*9���N�=x��X��4@�1�M�����*+h�O��#}�)lȈK�7\�?��g�� Rn~��Qڭ�aA��1��MuA	3�Q�����~����`q�������[��#[�}�`���������} B���H��,�ƀ���)�ؿ&9�;�G/�u��L7�����\0��e���yY~�|�˨\��ra~�ǐ W_���7o���	�m����}�ҙzǷ�ڵ�og�[;�I�]%����/������t����!K�T�Q}��i��C������?�\��@���\���;�몲��$�{n��q���\��
�M��1W�����h9���n���ɽu��~Ex������Q���Ff'A~�u'�1��~#���".�����<?��j�{y^���t�_�w�����U�E��2 �U�}�<6��[�j[�!?>#�3�����֟����\��"�Z��Y<]S��RD�
�i�t	��wCo�iQD`��/[�0�Ѥ�g�Ίm�i Pd~�"Hj����E��C	Pj
����t_��È�~�M�At���׿�m�e���;�����n�����e��^���}�����5����i?���~c^?��������o| {⊋�-�(�P�B
�iB�䔾����7���+ܳ���}���C�IM�s��6�e%� 
@ c1����$�<������� (��DH��:*��ϔ�Y�W!û��	"��&>?��Չ��<
���o�d��]j��a�<8���SM=�>gy�6����Uy�{t��""�F#"w��W������_�8a�9�K�������Iڤ��1����ݳݫi�'�SSxLS'e6�`Mw"*r2��a�����J+�r4a�\���1`X�
((YK�-I�V��g��@֋2.L$��{�y�%�#g����$���Ye� P�೟*��?F�=�N0(���b��4V�Y��$$�Ws[1C]�h����,١�{ `�"3i�H��B6"ԕ�320��;T����XV	JR`Ll�	�zgJL���K����S+ 5\�=A�``�����G�KL�^f�s̺v��C^d��V%Fl��k�z~�����b�>�&��lט���O���ܟ���m���Fm�Y�;z��~�{Q�b����M\pK	����e�c�y^iQ�UJ�&���@E*�E�G1rQw�j�MG̱*o���T�rs�PŘ�1EO�L�7�l�D�c�f�����I_)�����q~����4�85��*��b��J~-,��4�$�,��?�%+��{X8aN`��d,P��K���.(y[���Y;��Vl�o6��&Z��rmL 5��9L���(��/�bP!,�ć��\|}JD)�^�w2W�Vt��(l��b�T1�J\kƖ�ع��3^��P��aP+	�;�K�G��SJ
�G��7�d�CA@���� ����Iˋ���F��@���b�m
�Db�B'�ԑ��F���l7I#S`ͧ �͘Z6�6�Q�'� ٴ��u�5�Hhnsa̢ڲ���0O7�F'����@p���t��y����:&�����]s���?@�K3�l7Ը������L�ω�i? ͇���kn�(��?}P����o�1����s�����`i��,��;°\������-܈���+��_-"����x��a���.�G���K[��R�n J����5r��.X� e�T�,�
�%))$� %>�Xݛd1�|[V�@j�c��
���o���#�٘K��i�d�������4��h��ъa���i���>��ƥhК41oxkS2�O=Ͻ�|�˾��a3�S{�텶��AI�/x��dW�̔aZd���.���	�l��?ߡ��?<��ooww����홙��1���uF����{ns��Po�f��B<�a��5\�,'�2���|����{�8�1|{��Xw
�J4�ғ�-:t�ӧ!
ճ4�M(dm���1S 2�M5�>|��>|��Y�������ps�����}�6��������8�����W��Z޸
��W�����*� *�^��:���@�k}�>�؞H�qw����l�@�QN�A{5���xP<��>p*�؁����� ?p=R�z�@��`Ɯ~��?������x�tǲ?�����~ F�W���O??�e��,5Ju��|;J;�����4ce����y0!vw���\�,�[��hG��w���l�G�l�*yF�oGx@��y�t�D~�<#�Q�/`�e�@�@���{�lv�E���8dR���)HJR���UW ��JW�������r�\^�_����ժ�!Gpx\.O���p�\͛pUJR����������_C�`��)H�k,8ׯ_�JS���Yg�����C~���e6�l���m�8���?�����b�f�	��i��ye�����a�!^����Y�~�ў������5�S"iQ��H�R)޽_�����������za��팟��������a�+� ��������!���u������(� �PPPPPPPPPPP00001�ppppq�c0x<,@��B�WWWWWWWWWWWWy�w��g���y���E]]]|���������3s�999999996&�儤��p{'�`X��X	E�`X�,UUUUU\�\W��������������������111111!���{#��s�;!����0͞�x^��QE�v�^P���!)�����/^��a �x^�/����s���w;���PTTQQQ<7���h���JIû�w���?��/�c�q�8��?;���n��w����П
4�%D:Mk��UEB���:@��t��:@��tE"sssssr�����߱��~?s���w<hj�R�� PR�� ��l ��l��.���.���.��x@ Zӎ8✻u��:�8㎺�N���T��}�y�����lllllAU4�M4�M-�O��?�����^�W�"f









	�������s���-��e��l����D�DBap�Ç8p��pi�b�{1r�/���r�g���������������S)��e2�L�S)��f(����Mi"���3��g��������z67����WW`k��M�_UBT��k��}}}}}}}}}}}}`�`����֯E�Lo�P"���k���aqx��k�����?!��~C��o���d2�C!���͛6l8}Ⱦ��۷nݻv���"}��`>��������������(	0�A0>��PJR����~?��_�|+Vߎ��������|���?���wffffffffffff����?�7ws��^��^;�x����y!�<���%�^��^��^��Y))))¤*B�*B�-!D��J��P����i���^���_W�ᆫ��iӤӧ7VL�ʢ��RSWU��'߂ A�y�.��꺮��k��}_W��}\?W�^�z�z�r�����Z�jըj��<�/�����|�_/���y��~~~l6^�O�������ա��>W��y^W��y^v�z�xAAA�f͘f͛6lپ)|R��nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�nV�n
�QQQQP**,.�[���K�V�Z�Z�hЙ2dɓ&\�g3��t�].�K���t�O6������`O���������E�d���:)H���\�������mX�R�~YEX5]�k�[�}�h���X��z�?���tS�p�.���&��;�/S�T�̥��������/�
S*gsq��=�_6�S�`c����.IrI�rK�\��$�%�.Ih���T%^�����������j4h��<�y�x<y�y��<�����]��>@;�wwx��3�љ���4n���h��}���l�h4�Mx���}�w�]�K�Qw�#IG��=�e�J%�\�='cq���l�\�**�ʸr���*�ʸr���*�ʸr���*�ʸr���*�ʸr���*�ʸr���*�ʸr���*�ʸr���ڸx�� x�� x�� % x�^/����x�^//����<�S�ӊqOK^2��F�Q���.�{�X^�e�P�I/"IL���H����<[���x����<[���x�	`�惥~X�b�,_�jբ�:C��q$�Hr�sT0���<���D��;ρ��m^ ��ڍ�ڍ�ڌ�y1�1�1�1�1�1��O���QꑨFZ����,,,%e%%l%�%�r��--,%����~~}}}}�%�bŋ�Ȫ��\5���z����׮��lX�bŋ�,���,X�{�d��"�7+�b��f͛6lٱbŁbŋ�/�_h�&��h��5���Ŋ��ׯ^�{ȱ<�y�X�T�)��T�a�B�*�r�P�]���D�}m��������m�����8�������q4�:�q��K�������>�����앾���߯������4��`j�^��?�:�롦�A�&��>7���~7������������s�ۢ��ݵػ�k���r��r�Ĺp\�t:�C���t:�w;���s���q�p�p��W�����B���P���[al0C.2�|�_/#&D��#��Hc�$�af%�]t���������o[���l%�իV�Z�jիU�z��؈�I{�y�^����,����q%ܠ�YbRIUP�����>�5V�f	��ä@,����o�����}������o����	�%�ZSL��OɈ �=SU5UU5SUW4uz�.�U�2dL�2d�,�,��,K,[�7���x�f�4&�	T��"!�!�"!�!�"!�7��D4�2	�d$�&I�L� �&��h���e�Zb)��Zf������|���D|��)����Gccc`��b�(��g&L���=�g��}�g��}�g��G���7���� ��9�33���
��0�Xf`a��)hSޞ����u�y#�
Z�)hRХ�L300����ִ
�j����A����~�@ׯK�)J^�	JR� �f�I���=�c��;Goo;X$��`�LI�I0^����`�LI�I0I&�L�T|��	��uTª��S
����v������awwUL+�?�L��Mq6�� 4�M5�͛.Y�f �E��(���
��*qb�� �A�3���i��5WL� ��%��j͛"d�^^�{�tL7���.\��� �@{�]T:��b��bZf@U%�p�8��C'��j�xX^U<�����V<����z�wm�)��W?4����l�I������aH�/1r��/���	�M��/,�Z=����Ἆ��.�O.
4F�~���Sg�a���ՌCl;H|��M��i"�o]],��(������)2(�n�6E<�{�j�ѢQ���?&�g�ձr^���v�y*_���/�rGq�*G�?#��Jm�#�����n ��\���5�W<�o��ۺJ�z�)G���⭧��Q5���z��nw<���]i�LC�k#�m	s�gy1ӎ9=޿�Ydt��7ؿ^~&1����r��4�~������u�}��>=��"�u�}�;"��A��2 �)A�D�%��,�%bV�0�!�:k0��%��X�&di��-���1�(��(�P�jU@�����W6���#���nٯJƲ�6ʻ-�a?���>M|sϯ���a�_����Ԑ~V��c-c#5��Wk�m
��)�����1t����k�K�������e�s_�x��5e,ir�ٵ�iT�	C��L꺺m�ͤ&g�����r.Sw�>L��	X\��.���t�5��,b�I�r��B�}�U��գkZ��w�&��L��ڵҙ�%{�b�Y��i�\�ԁ}�n�~�7o��v��3Ȁ�C�h9׶7�������gv�U�SK7���[�!𐼜ŃˬrF��6���q�S!�9�P"����5��o�9[�?+����wo�9I��h߿�P~��r[�azʐZ���$ECM-R�f2��e��b8���(�z�c6��6'A�Q���<����K��p���/�}�	�{����!,��)���g�0�l�׮���_qU0*5�pk��zX�N'�Մ��v�[��>���7]�ZB} sm�A�~��NZ^�I>�S��A���l��-Ɵj*�XQ��jV��o�}ש���x^x��DLPXA�il$l1t��Yg��t4�+[�v���Ms�R��˛g����ZL5���J0tML�A�E����|�d���[&fZ����G}\L레�LmvT��ddE��"��*s)F�ƳZ,��j��D��a,t����4�b^�[���ݲ�[�Fz�sy��,�Q\�����l�ih]�l%�+\��%)2�5�][j"���Zg�ok'�ũ����q�:�O�~����z�C�u��λ������J�
���}@k�O|J:�kb�O���߮�������'��M���WZE���v�R�W7H�I�B�;�Βb���I�4�כ'D�U��`���S?D�h(�6�X�:Le\����<��m��Y��(4�������/��D�g�-�����S��um/X� �{�OX@Y`��po�7z���"b�y�������mu֏4�-K�b-E��RS�d/�C30p��sY�&[�]:L��U߭�g�4T��o3�+��.�Z���v2��M-�������1n��Z�����ZvTn.�ݜ�ETP ��H���]���F�K�c��/P�J�j&u�F?4GlV�ϱ�{�v�Ӌ�Ƣ'q��BHu� �	0!T(f�@��R�;Q�a4�*н�](3��������S����g!q��/K=�_�.��W�ǚ�$ ܌��I�� ��d'������UM�U	FhJ��ɺ��!OA�A��.t�k�R���u=|��0/���� L�|θ|�v��4�O��x��;����E�9�]<�~��Ybo3,[�4�{����G^��uݯh���s����B�>xr�=b<Zs��p&��8�i=^/���續���}7 _�kG<�f�-�t+��ݽL�Ś���0^�圚��gz��03�j]-ð�ϡ��-~�����yǷ��S<3D���nE}�w��W����m�EnEX��K�w��ӵ�Z��~����F�{ɇ�}j��D���,��S��l͹V�Iك�]�+d�g?v��sbl��b�����2C>�mo���ǚ��cɽ�_����w0��ivM��mD��"��S�Ӛ��Z�m�v��P�-�yݾU��\�rF�|��w`�ȹ����-�.��փ ���>=j���J�]˙LLZ"�30�'���]}v�6uz�,�]n�sUW_���s����DY�5&����X��fc��6�բ��0h@@3T�
��k\�a`�rv�&���f��C^ޖSI��M�~��Q����r� ����Y��Đ��K$�^TZ��y�O=�������y����o��Xvu��s�?k�\Ώx�&
pg�\ ��f6*��k�-�9SXf�{�G���I:jd�w��i���(��6
_��A�3#|2ړ�� dGq �wm�-Z汘��K7�_����qw���?��j��bk�iX��s�@daym�b�wu��AV{n���o�u|��|o���m��e얄�o��;>ǵK����Yc�,o�Y�>o�����u^�O���J"no�K5�nե���%�����Vs��m{�j����n���O6�lסb�{҂�zdћ�^���{���.�_������(���]կ�n5.ioP�0=�dk��GL���]�݅���*�J�}�x^ج�春SO^�ɵr��Fk�C�����e_���gS:8�؏�4�3��}����20�[�3������2����ةO����n⹃ok`��?;����|nx���i&�eI�HHy�G�k+bҊrD�PT;/������������w��Mmz��`��m�$v#&4SKeo�4�o}�������}n�Q5�&�j�wi�Hwbx����fłc�P������Oy輧�i�5�j���FEؒ^��L�Q��Rl��o=���r������`%I5N�.��T�%�M]�swj�˝]M����q���K�Q���Pd��`=��L���\	<�UFp��V�*��O�#��,�\�>>��gOA�7�-H��֡�3�{eῇ&b�-4V���	2^������U��?��|�sٱ5JG1�730U(��y@ˋM�����#C������l��F���v�Qh��ݱ�r��I��~�������c�m4�M��]�Xٵ�?K����MF�<�c��682,�+`���l���^�|�q�S)�KN�j)=7���� юU ѡ�Ӹ9��r�������C��Y�X~�e�XOm���Y�����>�����r��5/����nd��9 0`K,�e��(�Ĳ�n�ןK�����vV�9�3���iߊ�#��h��fa{����2c��A���x��Ŝ��>M�7����ī%I=����Dq2,X���/JI�S� K�g�����͢>3d�D
���&F��^�жl��_�͙똃	�/3<1��bq�@ْ �㾬V�O�{��J��ܝ%�}V�P��j���m	��:��8�dD9�Ҹ�H �����B�Y&{
��t!.����@ ��,��d�&�6\�Hd�4,�Ɵ�
~���K�:���Ű#�X�2��>��a��Q]t����	L�A�z9��"�&A�o�f�=�/���o���u 6o&���܍��K���Hd�jdܰN���7���,���͍��_���{_���D��P�$��1�Z�;&FX&��R�����`��R����g�#Zլx��s�x<m��<��0�Ͼ���\n1��(=�8!�a��W�
�^����ꪶ�k85���x�Z�jիL�+w�����gh��'�}��b|^o��ߩ����RNd�)JTbB�O<��;lSH0 a���m@�}��}���`�D��+a���!�"�(���Y��N�@F@�!��Ͼ����0f	��?O 8 � b	?n�iv!0~�2�qGq���!��m��4 0ffD�y�ӎ8��"	�L�n���Z9��y#����}Ė0����~�V4Z�E����c�1���@�k�xR���������@�0b��I��ϊ����.�=��1|�Y�7���&O�M��%=���W���,C��X1Fz����}F8 �ǅ�	!�Q+Zw!��ce�ʻ�����fF8�דk���nA�d;�|tZ����Hz���8�{�l�-����zM3H�����M����~��0<�F�Qr&fуRڌ��(��
'�hx�t9�H�
kR��p=��t���6B�U>f��1o�l9�2u�D�)P�T'1Ȭ�'����ܹ�[��Qcǎ�<x���-��P���F���5˗$,���0�-�we���K�X�,�á<�<<<�Hzzw�/l�̮�w3mq��6lف@�3�q[6l'���6ʠ$�k�B���YP�s,������@6w���{�W���l���r���$ܸ��b.\�ƹ�z�^2#0`3�?����r�p��g��\�rڴ���;'ڱbŅ�Ȯ�
g>]"+V��h���|���_�}����,�a�̫�LZb�d��2Zb͖l�ŝ-1b� [�ܶ�-Am�T[rۖܯ*[R�����-�[���/)yK�[�֗�����y�Ӄ9K���x���������lT��is����@x=>I�8��K�Xt�R��h7y�Xu�=F4�PA|������p�0B=�d�k�;i{qE.�e���(y*Re3V5��X�k{�g�oP)�%EH؝�&)�/s[��`x�x�?�����|�]+��� ���C���C㇊(px��C��������8�"?��(%��ȭ�BK ����Hr�Ӓrrld��R�򒒎Q�����RT�P�8�A(%8g hRzА�3��"�{.�*�"&*+>l��f͟>Y�dɟ.\٠�f��cB򌔠�i �Y�|��f 32:�h�Dg`��f�t��9Q��L�F"��u�=2S�n���n����Z7h�����������t��_��C�kw�_�����ܺ~o?���Ig2A�ڄA��g� �!G�E3��+GJ�///////.�������~�����n�#��c�մ��6�v�������r�׋ki���M)mmmmmmmmmmmmmQm���<ݳ�R���m�R���%�!�!@�S�Q�Q�P<�b�G��P�?P	�@N8�@O��_�B����~P_���/�!�� �(/����@N|�@Nt�@%Dy>�/����|Wā�?>K�H����>��v��.��V��uY�fw;��s��s���[��g����n�<�U��Åcݭ�@x��bض-Bв-�����-iK)6l�v�E��l��J8c\�c�N�!���2���y/%�=�4�͠.yo�џ�����H�ϟԝ�����]�n�t_�fff��������66666,I�����=9Ahh�	�	�	�	�	�	�	�	�	�	�	}	�	�	�	�	�	���������1 b@ā:.�b ����lz=�i��͝���QU���R+-ZǫݳP?:` t�E�"z&�������>���>��40�6{+Zt޷H2>��˂�·�I$�I$�I�����m��G4�a4�佧i��^}D�H�$��9G��c���(���IfGh`К�@�(��(�r�>�$'��hE��E�C�B�M*^�N%<D��O<D��O<D��O<��~O����Xf��:|s���F�`��Ϟ,�K��N���A�4�̒���g���M4�LԦ�3"��i�)���C�뒟Y�L0�����QE8�?����
 ����U�>(�~���nz~�����~�/O���<�`�����;�0`b#pD� 8�e��o�t�U"(�ӾN�;��xN�;�M�/��'|��Φ	*"rz�i�����B���8�(ۃ��Fq\�g!��l,v�l>�m��m��g���v
dB�o�ښ���������������L��lļ̠��}���Իݮ�e2�L�R�q��i�`tu" fn$d$�RҼ%�5�}}\����}�1��x��x��~ER���P�(��3@#1�<�b��W�1]��\��p��P7�C�<�l�6�"�qĸ�8_�a�
���\�L`�'"��xHFzQ��A�叼;�p�0�(�����Ǯ=��a���q�@���x��?A����4Q��!�FHIIIII/�����+�;rd�9��ZZZZZZZZZZZZj�q�r�LA�R�r����pm ����50a�8���R�Yr�΃O9A.�9��H��2SL4�M=7To��IH�"����vS	��i�ni�����P0DdFJEb;&F��e�,����+�� #�F���`Gq�Q�nP#�������Gq��nLB@����-���X. �8�6�8�񑝸�ȳ���]u�?dL�:\�|� ���+�!�t���H=4f^z��M����O׳|'q����ӧgf���n���`z����׭����Q�����ҝ�w����h3$6?�SP%��?N& e�ډ�L�8B%}��0�d � ~dBa׃���ac+q8eQE�(V�� ��u�]u׀0fnF`8ˎ�q�l6`����:뤵-anTfRː���l����8L��` ���)�����WP7����:�;�e�W����@����C6`�YC?�>}�˔1puB��ߦ�q5a�+Є3J�U��@�����gs��!�f���	�	Ff��6����9y<�VMd�`K)w�2�	'���Sۼ��<�#�yO)�<��ᰞ[_a��1a�^�у��-�`��)&+�WJn]�~�������:�����������D�!�Og5=��a�2{9���(�糟#��R&2C�q1�?>���?|��e���$p{���,�m���8w�pLא,�o�� ��01֣Ե�ut�wY�	O�|�	{���O&L��/�}�a�!�e�+�T�xlτ�gI�%�	�MDfYI^a�)��e*�� ,Az���K�ݫ��Y���ml��&-�����M�����)^41���Y�tj�X�^d��h�J�"�F������>�M��&�G,>��C��d�k�c�;;������ۓ�m1�o��t�_���j|Ki�g_7C1��p��i�G�F�dG���t�+���	���,0:�w��A���Q�sZ�Yqzo,��ù>7�m�y�S�zW��|��^셟6�'�zG����F��`A���h�̉�wνuӽ�c��.�>�3�9�3��} ���k�F��N1��CC�1�1�8��#��@��ZaM"C0�B�hb���`@�5�r|��y߭��liϠ�ƠҚ(�H	�Or���`n?����C��n�NKS��x�?X�����I�"Xa�5���H9b����[���x����MF'�2t������� ��A �#��À�AfDv$��z��mU�_XҚt�ӧNMy�L��5`����a�k��n鯯��������lW;(�����jm@$IB22��qA#�8�(|�}�L���DbeDSc1�$�	��8ɜ�&��M4�<�E;(�ƻPSnI mBBA/i����y�ѽ�;۴QZFZ�u���e�Hβ��W0��u�٠�HE&d@Β2Q�ݔ	�ifL� �fI�)�J��H&��%A�"H2m@�eM;;;;8bw�5�IEMn@�r������֥�!�!��4ȫD��0�:�1Ӧ{���O��`$��(��N,1*������=RI�J�`r�����T��7������1�t�&%:a�0�b(,B$O
^T���]۫f%
�QNQ���$�N9Qx�PFء+�n�C�I��m!�$�t�G*���n`�t.�
�4�|g�ttjmY �)z:'C���.�j����aJ�9m���'$��yqi��aXcL�fR��NHU#5k/��TF!Z��W��Mٽӄ��h@d�Y�l��"�-�[j8��sQa����@�B(�RD����E�%�c���s@� {��!ɜ	d��p��92����4�URr�+�=?7粲��������ݡr�U�j�fR�.ey���� ��D�I�!'3+�X틎�f���y�{�=΀��'2L�P�� $@A��F�"�MNt6�zdSV¨���ÿ!U�@A�Py��2�-7Tp�z7̍�uE��~z��%Ư������q^1TT�C�=>�{�	D!5M
�Eb��E���>�4�m�jPQ�V(Z�V�\�m�TX��
���Z5�� �T
���U��Uc�QJ�DRЬ�(��eR�R�"�Q%j�PDm�e�J��+���PPWF�X��m�1�e���n}��������z�`]��Q���_*O���Z���<Q�RW�@\`������x��c����Am0��w`4�8����+2���m6_|�����<hF����e����qn��Lթ�$Ƶ/B�w�X(��̴�.6��W��ߎ���Ql�����]�|Nz�	߰�  ��w/_~���	I��x��o�U�.g_ym��x����8Auq_�����:ׂ ���i���=O��@d"q2^���<)������2ݜ�gFox'�����$��{��z��|�������p���� ���'�H���_�֘f_�v�c�����e�����g�5}�d{���[�~�w�i=�OQ	u��-?��DA�>�Il����`�7_l��Ʒ�7���^`o�s9	6GU���%k��<86��b�X��}+���C0�������i��VvCD��A[̏��I�~�s�C� r�
�������YWƼ�z.G���率�l����`��������[���� =�7�Cp��z�ʌ����x��:�DAg\�z�����gg�1��@�LԐ�u(e,�~K�T���k;�T�t���v�w)L�O���[o���۔�|W=��!~�>�|x��}�Q������йދ|�F{lG�i-��vx~_ϹkB���u�^�ru��t��o&���\ױDX=غ�>潰�`�a�!�h)��+9Ұ�P��5����N{Ϝ�~HCc�-d�&��ܳ��fT����CŖ#ÉSg�E�#��^o�N������ܛr��F��c	�I�� �b��ڤ�{/�����ܝ�����4;�ez�Qz�s�������UPK�>G�z:��)s��jv�ZW������Y�\1�*��H<��V?�؂~݆ ���`���y�z����=����T�;�ٓ�򣃤��ޢ瀒�푐y2����*��M���r]k�v�MW?#�hr�a���>�;�m���"	��^ȃ�z)�#��E7��M"�VT:l��>��}P/1K�|��{�?�칱]��˾O��0����:"`��O%�T��cL�=�
�p��Jg������B��6�{����\�I�L���C�0� \s�F�D�u��<�e��z���'W�-���������*�x�u�vU-\�]����n��"!���$ �Ԁ�c:l<��g�Y�'���A_Õ�O�H���pppppppq}�'��9���?I�w�#ffw��
�O���}O�c��߃��찾��6L@@�Ҷ�Y���<6�5"�W��7Èq"�L�@�X�8ʌ������ύ(���A�z��
��Z3BDc���@�P7�v Ɓ� *= arc�th���(= 2�2� }�0��6�j_Q}��`�%|���~�������ߎ��a�A�Ī0j @ �v�#,[�՗�V��ЬKT[���XZ�Җ���4Y�2!`�_�Ͱ]�{�Nݻv}d&&L"��"�T��R*EL���w�w��y�w��y�w�坜u�������������������������������������['��d�V66666666666666669,�K%��d�Y,�C!��d2�C���a��l.`,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,p�&0��c�5���Op��]ˎ8�q�m��q�Y�q��Ok껿;���_�~����q����������:��s��3*���fff`�Ye�]��9f�Y�[[[[[[[[[[W�X[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[Qc��l>��6t�Jk�=ʚ�������l�W|�w;���s��~�؏a�ؿ���޿n������0`�������߿~��c�q�w�q�G����ַ�F�4hѣF�65���cխ����F��>v��ϟ>|��}��ϱ�>|���ϟ>|�ћ6l�>����џ6pz�h�3�ϟ>|�ug˫F��͛6m��ϫ>|���hѣF�AZ4f͛P͛6lٵf͙9�f�U�(͛6lڳ�ϟ>��mY��N|���խ���+ׯ]�r�˗�����h��xd��F�Q��j53�ɇ���!:�N���q)Yfl�T�����ܩ��]��m��/jf�0fffff{V�^��UUUQ��Z�}����UU�׳���˻�����������������������{�-�~�:NE�)txS�֢�"�'���}f���]ž���t�u>�g�H# O&�v4*ױw;]\��O�r�8�(�;��.���]���U�X�Y���Aj A ��K[�v�ۻV��{��||�_���Q��E�,��I z8����o/�ٳ�^	!� ;��b@��1����� �X���❯ĵ��XA�� Jb1S"�B�`�g�������@DD<��	�G��5����Q�Z��m�#���`� S*e�9��i���� ZL����[DX?�پM!�i����s'Ó�8l&�k��������B-�.-������J�Qdqfs�P`h\#p��)�ݖR'��z�>?,W����a��p�>�&/o���7!����_��r B
VVV(�eenr�0T3)bz�;��e�@ #�5Fq�s� vD� $�!�o���˰�Ѳ8)��l�����w�bR��:M��w����W���n�G^��ZT@�@?�,�~�ij݃��<�G��)���{��Z��&O��{�.o��OAXe������y|�U��k�a����-��gw�ы6�7��M韁�7Z۳%�/�.�X,��r{OaW�]�/����o6��;;�Q[�^��=�.,i��oܦ�dD�n��˛E���A��G,��kF�ǹ�Gw˰>|;v�Z�.�
�s^}���x Sq˱�fV���<|R/�!��������A�������R�z���!ث.�}�l�9�\��q�[��R�]粳M㭃o{F)c�ɷ0�ٿ�J�v����v�;���s>Cr�7 �C���y]�g��}�~H9�� ��6�Y�t�\N�nH�n� �T~}���	��(͵�l��q��z*� �� 840B!���Eg�:e���%�L� ��A�<ʁPA��$�؂ m�b�H�y[���Q��~��Ԓc�0J��=3W���W�7n�/;�_��i�}��4�y�<p���s~�ͷ�������z�'�7J|o�����o���l.���y
^�2��bX��y��Z�����걣�#E2Q]�njі���mľ�YCa+�e��6u��l/̵T�<ݤ���X�l���3ߟ��_E���oVp��Лk���u�̃:�J�Օ�4.�e���͚�e�շ�V�eݘy�9Fc��:�n���g��'���@�<����W@ѥHFrg�G�z� vgm�7���>������n����f�����#HD0*�� ~��ЪM�L��`<�"f@h�C��&S0����2&dQo�∡U�V�"E�Z�0�w�>�E��b�0`DL�0��D&n�q"eo)�I�,��q�[J�W�UV&!��G/�a���S�WD�ݳ�������&��}���_��>����>^�m�S~���<ӪuԺ�����t`��H\U&�"f���U!�=RzH3
(� G��z�kDZ`��]��x39��
9ü�hp��P,]�h*yg�V�| h�~�,��Y��]�a�8b��o3p�ϟ�9ˆ���a�;5�����#2�&WB��T>8�� UH�⪽2 �z�� �#��Uk����b�wC㋺j����To���q��x?B:t��n8C㋸`�R>���� ��b�UdU �5�ϐ����3
�2����wV��5TP��i��2��ހ�F��ʆ�.� �B����n����؄�}D�@|>�H�Y`�� ����%����?ǟ������.�*�U~
�v���oB�3�E�� `�n. pP��^<�`��kJ�@�C�p�ر�6.���,)�u"���C�k��zD��$
�pCcL�,�U�c7����«tH�֪A�gz�Bi��p���hJ�=��^��_=Y&.8�S!����5��d�=��_���}{�^�����]�0�mkٵ�.ܑ�{�񫺾�{����B������!�5�qrO�F�e�����8 �.j��w�Gl�|��Z�݋�a��5�����1�P������nph�9c��0f�m��tn���1�43@̻ �[0f�V�{���F���$v�`��ps���9 }o���ps��Ţ�6��陷�����8�Z0*�9�)��؊�-�o�.M�AZ6�:ޚ�/"ua�?BY�#����,y[G?��?��Y~�� ,1#ay���[EQ71,�J �9<.��?�y�|/Se�(�J(��>� �sB�o]���(��(��&��kƀ$�����0�^�@W�DF M�`��4�w9_:� @� Ϝ63㵵�	����SP/�֝NEɋ� q�@�8�� qf�n»π��hr�&d�N�� K�`��Կ%�,�/4r��8�&�hirn���G6y��s9�,.llZ M�
R�߿~����߿~�z�߿~�/߿~��N[$)�f�}� w6���Ȟ����ۻ�,�݀a�ھ���`5��0�n���������P{�����c�Aa����J�����e~D�o)�����u �)W*�1<L��6���pू*��E��:���",� ��;/�b��p�;V0�	�R��/W0:0�8� �0P�*���":�q��ᆒP��@��X8�q���N�f�(-
�)3Ry���0#�0>�) ~W_�~��������w p�25��6�m��n `~����������0�� )~�C�{�4p:�$�I$`2��g�f����<�?c����M�px�MM4�i�j��bZ�0:�>��A �O���<��>��D |� !dC0��A0�� u�q�H6apï!HX�`&$r��u���H�C�^�R��ٮ�h<{0%�&	�`2�� �we�ݞ���p�P�E��b���R�)�t�p�*��x�y��R\L���ai|�paXN��1�J0*Q�9�i43O��Q���R�+;�Yɚ� ��!�E������ڔ_�P,߼�������p�z�8A�o��7�����7Rև$wN(���A�|���������t��/���l�:l��l�ʬ�ʬ�ҷ���6l������� ��`��&�i������Xɴ�|��܌C*DD'X(�U�W��N��cs9V�8}=v�F�*�6�F#)p���LO�|��N��F�6/���ENǼ���t02`ę�"&�t�>4��J0
�I�s�|�� A����xp}���s���j��܊]ػ��X�[3fu�=�wF��H�&�ۡl4ޏ�ps�8M�"��e������ w�?�� ��� %������B�DJI�F	T,`,Uյ��Y�[mv�]��\���o,�"�a�����~�����L�Pp��R��9�M���4j�L2ϸt��f�Ba��d`xKǾvP�~����
�����}�f5� �H+�5��/�_�~��3g���P	���� ��K� �za�6��F7$9I�Q �����q��>������`f�����@T � ADA+@�|��/��^c�y����	Nr�t��y�V4g� �15b2�5Fq�jt��MQ��Ϡ/��Qư�8�f8�Hwy/����ʠ�,�$H�$�Ik����gd$.�E1L)T�D�YT%�Yel���0g	�Bp�a�C0���B	�2�*1�x�6Z���2{Շ����P����l��n �Ǟ��}�|���r�(��(�J���ŋ+EU���b"��2��Z���Ym��U��=�;������� ��]���Џ�)w׏ܻb|��/aR������;��:�a�����{�	��(7zȟS��q&`Q>y��sڌ�OͿ���6� �U����etrn��>>�2>6���"5��z���YG�v�� ����:��#�c����v�='���k�Y��n�ؿ\b�_��O��D2�=eW'�k���V^�J]��zO��r��������_�mz�[��������t_��uQm��TI6�͖V zf�ߏ�99�j�0��6���ea�*)S���Ǳ�����g���b�i�i�=�3A*��(1�����4�01�Sp�cޟ_8�Q��A�d�|7����ly���*�}������E˺��u)�ŧ��Mo�n;P�O�>K�x]����io�d$������ ���p�2�����(��P��f�h�E;�����ĈR�HI(���E�T Ȍ"�_�<g�|���IFK���>���/�
� ���|^Ӎ�������7?��{�'�m����˶DE��+���!��$���_��(�uG0uߏ��%�"�mr�ﮫ��/��ON���#r���i��Yu���K�z��UX,�dӉ}-���39{Χ�-7�Q|�g�۫��?��k��ù�`�fFvd�*�=5�Wԫ/�{�������&vZq���owb�6k3�i˪��|7��y�Ȟ��Ց�6~m�g�*�ӻ[^�ݗ6���� ��V���R���7x^���>��X�2#�wjJ�;z�g[z�Յm͆��c�a�<�g�P]�{.=j�i�b�����T�pk��Nw-���,��X�.��*�P��6�0_�Xσg��7����b�R6/�ɽ�{	�b��MMm�4��%�'���j��Ϭx++?+[M�pC\4ǭ�Z���\�h� $�F �� ��qwz)t�V����+{�gx��ִ��%v>�|��_luGa�R��q�+���5�R>�~��~��#�vїn�k�|��8�x�P�'V��m�2�5�Y������R�6,V�o�w4�4��k��0֗5�_]Z�8����k{�0	/7�w�ʾ�ȿ�]�QLiN����`�����4h_;L�����0�J!~7�6�m �+�o��n��kk0A�/T����hq�8�B�N9@�*��Z;8��`(�Z��E^,�T�(��T�UEb �UA�(��f	�YO=��BBň� 0�bz�X�z*R��"r�������/�2���QUD�`�ŝ�j�-�mBШ��B��ϸJ#k����Vbb��E@��C������H�;U�Lj����_!����܇,g��C�')�z�P(u�2��+�]@4�� ��}+����`�Vz��	��t9�^��>�p3>JK��aa����sxl��I݁��oXM C��V�S�'��N��Ǆ���@P�q$Y}P~i&���p9���p��C������d�j�b�{/�5�E��?���%��Wk�{P�?��U惷5h�O�`%��А�����p�ٳf�~<hO�a$���w���.����v�q��7�1���[�ʹeL�q��X*ņ�,lu��l17l���.ZLCy0*7�DK�2 �#e��~���^W���[1�,�V�;jT�F�m��K�����C�#��.��ڎ*�Vq?��Q�"{! K-�K@D[R�ԗ��+L�D����۾�0{u�9�V�%k?N�:���A�FK��n��<8��=R�],��d`�"D`W��%�?�ѳ���g�H�����:��x˯����wݻ��^��;�F������wo�,% �61�l�(Mݛ�oQ���nK�����%��>.�\�k�m�f�S�ak��Jx�YL�Z�q�jW��^��N+xl�}�暼kCŴ��w�)<����U����k���u����Y�Q�2�4.��lo�y�R�˭����E{�R8u�d�y/`�����ܭ�N�yW/�dȊl�Z��(�Y1���"I�O�Ӫ�ڵM3������<�"�m�af�|r������n�����ſÓ��]�sV���`�[��[j���%���ҮS�qe��c���˻�em�<�V5M��M]��^Y��/��Pm�Y�e����ｿ�ۿE�z�q���W���j'ױp�kZ7W�Ud�N�ߛ9�t�Q��,VCG�n�]�tc��l�-;�~�]��0���-|_"Si�V�����m�u�8�0/ץ,�g;y�m����ޓ6h��]��J~f^���7���x����̥��j��&�y��6='>������f�5ͤM�M��5�w��mMNh|�1 �H�k��AK9Ƚ�DOQ�<x��*�FE_'���*�2�� t�_鋁 ��ԡ�H���^�ߟm�/��g�'���K���PN验m%H���	_��1�?�s%E�3���Q?x�dA�� ߻� �k:.7b���p���E(��8�Ffv���S�j���c�&�h�@k�����z~u������������!hD7V$C�fD1�C	�"���g���i�2��Ђ� ���v��a�z#���7��%�EW`��Q��"���|UE*7���Q\�5=�m�#�>�.`��\���/���B�(U	Q!�r_��O����s���<^o�l�����G��)\"�W=*Ҫ�|�	�o���>�8BA�J� y1� �R��8����]��4��y����P��������ja��<g�4���I������]U����:Z�����l�i�ok�VGq���K��2��m�mk|(�!�����+ў�|�Nw-�f��-V�J=���n�m�#R�X�i�7'=�p]_�[��V�f+w���֟/��)ܿ���ױ���B��$�|L�:+�qϲۺ�&=Cl�f۳��j�2f=���o�^]X!ѫ�f,�ܳ��ߢ��o���ҭ�t1�Oa��M��cgV��M�oj�j�M�3��w#5;���찳{u��ݎy)ШD��o=6��ro5��~I�{b��v�`����5��}�<�wn->�>'�筚���=ȫ'��3?�wyL+D:+=j�oM��[x*����ۧ.������i�jU��G����<y�8�U�w5=ǱgbL����-nE��಴ܞ.X�� +PE�Ck0�U5��k�פ�MU�-��~�m����ln��*&_^��mɪ����>�f��&R����Y'M���0s�6o���a�6��e�ڼ(���J����"�㵈a�n���,��׽u(;������$�Yı�%�|;��6پ�F��䎹�d���}�_��q��q54kr��d�����5��QP�F	ݜo�a?R(a�����{�`/��@�_������h(�Ŗ�(���c�PX�>��0�Yb�,R��l�F�̳#(�F�RҠ������~�_�_+���~������
vG'���}Ao�(���.�}�Cy]��V�y����$�pD/Aȓ���c8�L�#ͩ�����)�)ܩ�����
p)����S�{�7������b���(:��K�X:�ȉ��>YU�2��G,��R�����5��^�.DX��v�~kg��V��6Oz�.Wњ�|Y��ŗ#p��~��$�Ԁ@̀/l8[Ye����*�.b������_�����`� �t�W�;��hYr]�f�Rɏ׈���<�.Vn"8���3p�y:�ȁB��C��L<�	�l�Z�$EMpYfs[_!.ro#�<����	�t�d������;ʍ�
*���aЏ��)�<F������)g%dB!p��t!	qb��H��
 ��G��K�SN�m�аhYت]N)k�l6��Q�V�������}Ș��2^߆Ջ�9�g�Qg�3V+��1_�{�mnA[ۧ��L5W������n{���`���.�R�<w�M乯8S:d�o�{jlb�ּ*b�v�����K����dj����Y����lNޔV�ul���;���n?s��^7v��^�ax7`��g��]5���9�墙z������0��iaJ��|T�i�y�%�۷�]�v6w���M����u����Ɩ��j��Ӈ>�tc�ޢ֝�Qw��,�L��7.n�F{�'{Z�i���9.țO�+Y���|+�].�ݬMږ+n�f��+���9��~˙h_�B�TJ�Ni�_.�m�W����&�\�Z7c��M�{��!�-���n�i���Si�;���8~�ܠQ���G��}�5���sazŤ2Z�M>�V:�MC�f���m��r�ڦ,\TUs���gZ���xƎ�Oq��C���r�õq��'h�ݧ-ӅW��6�a��b�L"�
��Z���hi�ʬ�wټu���^5�]��d7,@ѽ�ycZ�bq���y]�N����߸_����������$�I����k̊qP�ڦe�1E��e�-Z�t��7NVϯk�P�A��`�F|����蜇\��ݜ�~�~8
�ǔɏ����c�����[��)���W�w�W1��*yu+ѩ����}<9J}�eNR�MO�����1N���dS���*"�x�yh��z�=��:h�'G�p!��e@ռ7����x�⇸�����P��|�<r,�ujɭ�.L����ѭ�<�ȶ|���i �I�$@~%O��?G�m;�0@�?#�~v��N4I	2B%�E'ȉ�{���������v�7fp��2�����<�F��b����~r\l�p�UsXꪣb���}ڑ|�P����j�k�������x��4�����o.f�;ec�ʞQ��9/z�;YʮNl^����$�l��D����d�Q��%s�U�Lّ�X�8��l"�y�o���W�~��Q�?���~w�q�/W�Ng�U_�]T���K�e��!������P��`Q�� 0CWn��Ti35�9�	��Xc��`��n��3/Z����S��u�Ǉ�lx^5^�X��Vj>��$����XZ�|�8+�e.I���������OS���Q}u{J���ד/��Fn�푵շ���lڏ�dC>�n�z�Yk�=]~�����tT`��������{NŹ��-��w$^E�r>���u|ZuG��+���S��cl�vYp��{7��m^n��7o�iثO�3�ho�ߵvh��j�;O~�K׼�+���f-n.:�KS6��i��Y:ָ�{z���ۯ{Z�6�ۿ;[�̶ֲ\�+G�2U3K���,��<�b}�B�mV��J�kңoo_�i�U�Y{#ڸ�m]˦;���Ӈ�������u:ˋ<;q/�G��~ͻ�ͱ_u�������޿w�����ӏ�@u=Ϫ	~LRm�-�r���w���n�׍Kx�̲����y ,��ʲ�a��Y��~���]kv����i�iof�<���_`Qd�ط٤�Un�:�M��r㶚��y���)i��3LT]���c���I���
Z�uH�{��lΝs��m�m�Vf/���?|�o;K��<�E�~!�\��〬<�V�DJԊ�*��0\�32323G���r;�ߢ����ޖg���v"?���"dC��u\���w]y��`1xJ�!�����fN8�ھ������ ���,Ii=��eGE��r�a*�Ff�j���0H�yn�r�������0��y���Ϯ���iP�!I~��� �����dˤ���>
�/o�|}�2'��\5�.y�)<r6��Q_i� {>�iF\��3CI4  [:y������eyZK*Ãu��]�8�B̥�P��Օ�a�{�S�;�W�\ߋ���/Y�|�a��V�e")HLz���-��~m|����=\4�ʺJD.�"E~mv�M�@������,��/�,EI ��F���[���ZE��W��g�.�T~��V�{���f�IŊL=�۶[��k�۸�&l~�Z8�7,5��{�i�|j�d����7��b����f��R�5�4h��,�o�;���N�NllUs%�3�;���C��V�Z�u��6��/9��i�F�X�@k;�"�����)Yp��siʘ��kow,���+�������a��skL�]����v�f��֝�N���3*w���ɷ�s�~�x�����Kڷ��V�q����@�̓ږ����g���ů���Nmi�&󬹦�Yx�pZ�����kPZ�;e٭��"����\�O� q�A2#�h3�%��T�fUYI���,��(#>ݝrt)Qk�&��<&�| �����`�6���/ETλ��-=_����,�aVC3;*�!m���*K	��R��3:ѱiy�i
i��i��+Ju6�jl�E�*9��ݏ�Aw�4G`HH���j	Fj�=�����y��_���_�T����ܡ�������&{dߪ����6��J��R+��J�~���r�|�����w�g�z~'�}��w���	|n�Ҥ�^�UԈy�dC/��H��e�2}Q��k�!abB��.S�B�` F�@�0�X�J��׃�;<�嬷�$���I���a��)��}���7i�mk!"��(��k��7����݃- |���?���s�;z������^F
�������!�R�\�
�nra\�R��3w[o;R��JiT�6c�I^�����N��Di�'��w���3���������O�y˙�*��|��yt�]�/��0�����80�̮�I��͍ʾ�6��m��ӻ�;cy��Qk5�p�����T�q�7��v�ƾmD�V^������+��R�����ӼKv�9˗��cd��yd�>F��*��%o'ryZ`B5�$dZ��nj����I'�E�./���w�'6�g�r�|%hD���9�9��1�䬛�U
x^y��w<��j�C�w#��r�CªF�s����:2�oJ�B/�ޔ�V�-¯��2^-Bk8�q�	e�n=Dp�n�y���f��r�{���9c�O��f�̍�;���`��Q|���fFr#5뎨IǸp���#��������k����Z�'of���g���D���T��
c(iy9�KLp[�;ۑ��9y��>�Ӑ?9r(o*.T�3��S�/&T���Ÿv����\��ӽ�Fr��~��eD��<՚��!9p��K���|�������'�.��:�rDޛV��8�U��ˋ8�7g�6�����sg��1��Ҡ��93!qq�\艼�TL�J�-�5Q˥8����Q"��n���ds������?��י�rV���w�̚ɸ{�x�x��^�gN�|Xmٌ̜�_���8�VP�:'�a)0�2�X�O	}5W�Z^���sw6�M8�~%���j��	D�L~t��rQOΗ�=L���]�=:��gE]"㒬�s�xo���h8ѥir�c6q��̞���w����ΒkgD��.I~g9����[���-Kݘ�r��k�bO3����{���{yF〈u��}��̳Ge�\�Q�E�p�U;u���ش����
.��>�U^]�y��i�3Q��5vzoMˎ���:D^��Ft�Wh�W+"���pQ�.Lr��k��z���*�n5͢a�7�.A44�µd��[��(�.Ua��|�m���~sy���pfƾO,�o���"��yx#�o#���)�c������FB���P�w{���1\�Ȃ��j�f�'&�u���w�b���z�<V��f�s��H�qp���H��/���1�jv��N��n�b��������Ç��ɮi��'�<E�0�"Lrk��6*V�{O���\ܪԭ޸_��i��s_+wvE>�n�~s7��j�<�[k$1�6*�qR���/EM��2��4o6\�U�0#�̹�/��S���7I��e%gc��f@����n�����|�ȳ0o��*蓱9�ˋ]��;K`�{x6�I�6��sB*��O*����v��#���6����ҵqʓ����Ӄq�i�C"_��iG$VY:�fʞJ�{c�燊]�(�/ٹ��c������;�M�����l��7U'k�͍�-nE�*&e5q�r9�jO4I���mJ˩���Mo�UTn�Ës���炗L	������*
��az�,n�]k٪�B��⼺\U�B09BĎO�!FY	f���8d�]e)uo�Z����G$����dQ��m��6DP�[S��8���ڬ�4�dGN��+�|�iž���O<y��<F�4�n=Wb�)<zؐfvyy�w���_#[�1U�+5���_*c�"���T���u��8*.䚈��ʁa��%Mל����M\�lC��r��O3(��s ������õ��Ҹ�w8�A�GLu�k1��tpp������k�A�J���_��Ni�'�e �+//m�`����wy�q���t��.�prn!�{�Y
q�nr*�-��rfi@:��į9���K⨳3�N9K]�7��pn�*n�Z���7DP��w��.��ШD	Y��Qi�}ბ��=��%f4��ͼ�+�m��m�̸�Q����htq���s6��sc�nҬ�5Us����۩���S�Ї(C�+���;�@P�M�e��9��q�;.�9|;�r�ʲ8j�c����\y�c7t��M�7+#"�l���n�3��$=���	yڕUs�KU�Wtb�����r�2�J�	�*���Z�ś��0�q��we�kb+NK��i��r"�#n�·<\Ѻ�����f��0a�7ޏ�"�3�F#i�ERYDeR������]��C]���(wl����W\VJ�4x�}1����5�Gfn�XG%ب�7��og�^�x}�=S V��{��n��x�3o���0S��z������o@�����o sY�U�῏�����w8f����I�Uĉ��>���;�.˻�8�����"+�IF��<Z"�V��6�c0-�������x0ʪ�q�U͍���r��ZW'��2�͋v��O���V�{���7r?EqFmN�<�Tz���¬��m�NU��v�������[@����`ӆ+�5�7���t�1�O\�Qǟ^������U�u�1oODژN���i���U����]M�ӫRgi���o�N��Z��Ɇ�ue�U��L686krl�Z�ǵ�U��rqɝ�܊��l���=ʍ����_m�ni�j�J��k~��f��Z�F����v}�\<9dA\����z�|�F��O�^!�l�^�n�]c]g��2�:� A?�]�
�5����+Ҷ�lu�H����*��B�J����5�6ى�)�4�*�t�s�SKN�N4��UYT����u(!��W@bwLG46�H�Ȟ>	�H���@4�|R5�� {i>�z�����/s�t{=���:xj(��ƴ����+�8Wa�#� ���H'���D�P=�<�	�b������+�P�tJt]��<��v}���m��Jz���#�����e���#�
�@X�_�?%�ujV�$�_��>md��ZQ$�U��iCq���$][��B�ƄL cr@�S�O�oZ��)�'!��JC,�X4'��h�?;��]��8�Qt����QCN!*x���"���VC@�@��Y*,V� �+ *@*IY*T�C ¢��J�E�)`HJ� �6���⥢+""�E���`b@a ,	ZʂTD$P�U��D�d@�X�C���IP	XF��R,X) �� �H$XC,�����YR�VJ����RPdY,Y����PY"�����$U��x��H� 70����aJ�=;p֪U�&VA�L�Q]�l6Z�Ia�!��Tdq���f,0ǈFB�d�5-30+;�5Ŷh����Y�I�,�0ir�9_��YW)"�V�ro\�%�㲊:�ޗ��N���՞����{_~��=s�[������k���
��m��s��v=�o�q*qķ�����S��S���vs�L{���}��Uf鴱�5u�����ٯ�@�������ݹÀG�9���ǯ�{{O%����˜�	�>��76��f��s�y��=\t�����;xX��kG�{T���-g�n�� ����=��EF<ذWo"���q`��Ty�{�ݭ�:6�S��{C^�sw����µ���ɞZ����ɸoj�Hڬ��e]�ڱW(C՗G�q�Ǒ��srt[����[wG�&��e̲C�ʿǒ��Zݛ�36�<��|5�ۆ�<
�q�Y9�KZK�������C�.�}68��js9�9��m���9`��H��fK���d�*ZX�8�
S�5�Wr�}b(ь;qC�E�"�r��t�C` �@��7�����D;�gm���g��u}����4J#��� *8Y� �>���"]?E�i>��H'D@յT��X� �NЊ�n��=���P��Щ�?=1��i񶉇��k�!�����y�`�s���E淧�|"ut�|~0�|��<����R����x�AO����(Q'�!"���R���N�P�^1���2���+���[;�9s�����NEZk�����Ҩ�� �#��A|�T�J��F黓o���e �	���X��U���K��셆~���A�b;��

��&b,�c��OO淡cJ����h��v�e���[�4Sϴ�*#3c�t�6�:����~%$F�c��WY� �$º�`�|N!���W#� ����"' �E8� ��@�� ���fBOL��*���Z��g�w�x+{���>���iTU��~)��1U�?�����KA���~2��"~���xs�O�HD%��2|�F@́�n�*D�/V��{#)h6�l@���L�\�8���Z�m��W������B�;͵��R�5�ZcY���/������yn� �����
�+V� ����K|������"B�����PČHґ(D"@><u��.۵�2�?ϿԽ������]�u=���~����R�v7N�;c֍|1˒��ӫ�VM%�je���j�)���B;-E$�FA�/�(u������}J~����E8G���8���=N�wn�{���SD���*�^2��|?�av�6��>�h[��ͫ�o�$f6�)o��"Li�'�(�"�1@uB���$�i#���>S��ӳ��M��{0�؆�s��o���g��!����a@r^���O�����$9���F�R
�*���,!����ʺ�ϲ<�~һ"iJ�X�G�ʼy�Vp9��h�v������`���a�=��`�����^�{���i�{�ՉFU>��j>|.��9:%��_��3L��9���s =N����ٗ����5h�=c'òI߰�1b�0/Fj! ^O`��1�������S���K��������k/�v���=n[�������o�ɨ���7gÀ��PHtE���1L`�������B�AI�k����ߧ���M�Ʀ�� �Я������T�4 t̄ۊIR����24:���Γe��򭛑��30`\���#�<����=`�&/���ǠO�����z�C�� !점�j*2x�������[��U�k������N�t&��|S��,�s�y�~@M� �, �����m�j�G���|��:��s[�NE榋��?�d�Jr٠�aIT|��~��}���gn;�Bg������Æ�	3��5&�YF{��å0�d��a334�'>3 �$
�s:Ab�	-�8e����Nl��˛!�6q��o�Ƞ�8��L�!�A9��4	�d�q��1����ME
�7͆C��9�mb1FS����WZs&�̥LӘ/[��W��¸��;L��7vkY�n�5tuw�D�]�,���4�T�6&;]�y���)�r�/��t��-����x�Q�8޴l�D&{���ҤXvy,M&t\�.&.���+-�5�`hK�N"��0���������kNNoI��p�}�x����Jq��IQ5j�c^���ᮝj[�bꆍQJ�\1-��a�0s-r�y�5��f.�9Zp5sy1x�U�x���r�a� �Q9���*�*hvE� ���gf��j^MÖb�W]Ю�ƳY�f!8S���"%��
RPp���P��)I�Ʌ��xH;"Z:�ē)Eȇ��H�i�=y��G��[���g�p�t��s]'-.p���q.& �PTA���LA\��n��۹�.	��r�c �%8t?��{��K�kZӮ���˥�N�A��m��9K=t��䀄r.�v�ai*��8��Lp�ƴ<�p��Wf��[m9~#�û�n�N�רrET(�D����'h(bA-n��).H3�2���"I.|�(�A��_kKӑG!���76"J�9��@=�����L��oR�Cc�XI" �k=���B�(9����I�L ���1���`�ڪ�2������T�3��H;��)-p"'��E �P�|(� H"=G�y�kAl��ư٠Mqѽ��Km���G�
a��rK��"
�P���Q)pK���!e�D'���v%D�f"�С��2M0ǍSC�a����M"�]oZ@�l����db&�(\l�(kA�֨a��T�Y�SOFXg�͋V�64dg�55��V�P���Q T��0.:<�HXL��kgqD8!��Bh1M (�2#Fq�&4Q�4d7�Xn�3(bT��p�XQ��q�]�7O&��S�l,)4q��MaaK,-���	wJ�tXZR�Njk��x�6��-8�ް*MƤ�/�ܥ^�\��ӽ""j����a�3(�ff�Ř�"
���(�k+��2͚2�YZ#�U�z���C��r�[���F뫚�U`��QEzO:N$=Hh(;�1�b�T٧w���rڶ�Nq�Z�]iW2bdަ�:q���p�ir�U��;�NXn�h���up6���\�MZ�n+\q�2�p���;�s8ɸ��1.�U@��2�HH$�r �oMJ^�̑e�0��QP�@&�e<�w;t�s69B�w�4�2�:�m5m5� //��F�%98��)�����s@t��w/1)�P�D��sS1��j�D�5N��� ��ÂFRBD�$Lp�����='H�S� �1�������$VЪ2	���qX��M�$�WZ�FD�j�@�'�*���C���2�;�~����Q0��I��0K��B
j"�̗�.V��s��[h�%+�fQ�3"

C�I:��0�?lǦ%���\�� �{.��.����[.��˨%�!z�]Z�S&��sy[Z�֌�Q�J`�� ��#���P�3$����2��$'��$���l[+.�
�D �à��e��I��tV��')����]n7�dʈ�
PL	UuCҬ8�B���wQOd�@�f�p�`4!%�Z�LM^�.�vk�tH."L� D�����#Ɣ]DB�ɈZ���]�&%<�Q��V!A�� %� $�vw7 KQ$�8�ņ���%ǖL�I����q�{��VlIi�|��	:0�'e�Nz&����m"vчlP}L���>k���C�f��|�t��6�
�W��\�LKBS	��dP2D`���,`E�tt�D��Iv���h-�a�-\�3Ȳ��+�#o��c	<�c�~Y�Q�) �}�}����%Q�v��(���������hRmx��8^O���"g��U��#�`�X��H�2��>^� v����_R���>ӹ���vN�i��C�P"����^/�B�I�9��2M�@�`�ЙI&�d�)b�Z�|KZ�x�%��]JHG�����@���u]�=��6\���?��<p�ڲc�Wɷ��v�6�"B	.�HN��-h�$�!�+�'Ht<ǜ�_3��\�n�j��*~�[�����{�YzB	��=4@����XT �1��n�T��'Q��W�7h�hgB^^^�t#32�5j�ΩjE}�<r�4䘡圼�f�.5�,�w����k�q�Gϱ�!����)v�O<�|�P?~u�	��lN��'�C�"�=/��� � m����i>�������}��Sͩ�=c�O��Dw��^	�p�0B�U,@ķ��������ݾ0iu���t�S�w�G��=BWQ^��TC���4h����%�!��(XE��?;W�5�jm+����OCċ�Cԇ��(��Į�b���W>1��2��e?����T���ϱ���^�
w^��)=dmi�0\��ԧ�;��'q�w��w7wzCF�6h�!�X��d$W<�:::s�ր� _�̃�;�&a��;R�
���%���@>���)A�?��`���fQ� 3�t�Y����ik�*�;��`����b�T���>�{��E	LCO��HaRTG�%HN��4����`�螂�t����j�7���<=Up�pѠѩ�&�ʅ�rSH�$B5A�
V�A���Z��8�@v�oe*�>�k���( }��d�;����h�X�������Tr��Zt��6�H�������>�{N�gg��>���[�'��➈���[��ӱc,Qަ���D
Z�5\�s}������y�սU����:�>R�����t+Z�مI�:�ߎ���__���ߟ�׊�	����$j wP�~8�=F�U���޷�:U�ޕ�9��t�3�eXt�d�H#��B��t��{��,�hR���{*���]�O���)�w��K����h��r�+x�އ�`=��~��YMU���$2¥�1�{�_������`�G@P�f����u:<��3	1��-���	�E`���Ѡ�d�l�/����I��0<�w\����)�(�Ǣ���щ${5����ep�H12�@(�p�T	������7���B#�4Ν(��9��S_
�8�SBE�x�P���"������wYc1��=�B�p�nt�5��J�T�����bi%��{g�p��-�~���M�'�p?+������"5D+b�J��?��|O���$��4�iih�h� �EO����J�`�ٷ����w��?�w��}�������D}� P  2.I�{>]N��r������4EL�m*4C������������ӑ˟��p����(���ث�A��j�	D�	�@�����n̠p��`D�� Pɨ��d�MKQ��.�2hx�(!�[�]q�q�� �V�?�f�� oG�S�����輯3��J���H��G��ӛZ��?g�W_��<�R�z�\�&�zP���\z��c
y(%��G��0��
�,��ab�HV>����k�^�Gx���A(� ��3R3�Rj�-������>�|�p/`>d,��5��G�~��:����������1-|d��H$����N2��������?=[I�LB \������JA�!#"�)"zV
w�SZM�C�!�RD@l��O�@��"CJ�����u�o��5���~�l'���q��}�x2����ܟ����3L�5��~����ԕ�+�D�3C��G������71̜S,���~&6�(P2����ǁZ�^՚jiIC(�4�c�'�ϫv\����!g�r1đ�Ĩ�0�"B��<^iؔ0E>{8���|��v2�#�������=+�dc�[��2�/m
g8��qI�&��4�#ĲZ�T��N��u<n6=�����3������^c�m'��1�?JC����sr�%j)�Bw�g�OS�R�-�:�N0����8]F��`7�v�1(�F�I�=��-A�@@�b	Š�

�}t�S�G��L�p�|�2D��[-��~�~F�1��_;��,b8�D�B@���h��%�������i2C��D�DB��F��zkV��j�*�@�����%�/M`�	O�֡ _A���H�*E��Z�"��>p�
�����q`�&�2)O��Z]h�D=0:�	Ӌ��4��w^��J�J�ӳ��=��Y7@�|�y�5��C���7��g29�B e�����"G?�! B�<�r�^�
��e�qM p�_2�E�=t��9��s(߇�������a#��O��j.O�3��0�2���%)� @~(��m�hH.�b�m��(* fP9����Q�a�s^�7�ª�cz�7�p��R�iM��nR��dֆEPP`�(�K !	�N2���t�b�qST�R��m�[M��<t`mP��gT]��ǥѴ�P!�`Dw��f� ԁV�]�����3 �":w�A�U5�Bq$�k��S�|u��-Z�W@�֜k0uN28���qK�ҧ�U�.�IX��,(����
�6�B�++h�imTU��i�J�O8P�� Q�sv�{į;�V�N8���[J�M=�++B�Vw
��$mi©�3*��������3Ѐz�=uߠ��*�}�CĒ��!;=��d�ռ\�e�Ǚ��������-�O��YS��)�WwN���ש�M*�r�r#U�{�/��|ʧk�:<m��tN,ɑd[�yVf��VY87 B�N���� p߰f v�2o#��N6�m�oA�L�"0����-R���0���[�@��r�_��(߂����[ܞ2��hS�)�0��I�>�e�"v�u6���O1��Bq�ݡ��ۼ�~�z�Ū��ZY�(L��@�30H�T҃ō��"8�#x�b�T.K�.�Q��@���T�� �@lg������p��!'��P9ld�K�;�, ��a'��vY(� �[-J�G���o�o��?@��r'��������vëUv}��Vu6���̖g�"=AR/A�Hyf=-�!Ǣ�kGX�v8㯭��hC��B*Dd>fw4�,�B�$NLɄ���
ϋP�
�~m��l朰����ӥ(���I�q�lՕ�����d�A��x��ӳ��W�!0��B�UUB��@`��XR�A}� ������}�O{C��j��o���q/�)<AO�_߰%D����R��[�,g4��o��
=4u#i#��̶�V5HSB C�v�>����#��x���pq�~��$$B�A6p�v^G�{@9�!�p@���N%7���ȟ��w��wN׀�(�
��d
�)�Y�
 �rC\0������2K3��{��y�@�p0�~���}�0�h����v�������}zE��HR�=t w�gT�d�X��X�N���"M�� p�.��~��*�C����W���ap� -�y���:nx}�x�@�!�"܊���fԹ���G?��8�?k�R<�5O8H����E6��B� � �Ͳ��jP�.��׽�A,)��@����˷� *`���>u����J����!A�N��wo�ez��cU6��!�ݨ�Np�;z�3���l���9#�.jaH)$HAc������/��!zJi��91��cy�]�������2z��=��:J|��W򷇘���A���5��?�{}O������|i��d��S[��'O���>���A9�dTz�ΊB�+��B��+��貴B�@H��0�2�/m�%��!��0+�������E����z���Em���\����P�O��4�Pu�B� `�=�ŝ����Cϐ������[�@dd>_���R08������>'S5�44� */����
�
>�|��њ�ս�����i�:[~����~O�m3}�����ޛ H�Ǔ�}eKr	P閕�Ì������Px�	DP���6N�%���(�R�D- �X,Af�R"w�A�N2�\\�G��ߏ��;k���U�~T�����JL�WN��0]M,)� '�?Tl2}M�*��>����L�6 �)�c�XP��Dp;Ԕ�k�_Z_�2d���V_CB F�TY`��1dcL�%.�1� ȧ��O�ḙ��8���jȁ� �!`�o�?f��S�s`�i�$<+Kcj�*�(��Y%�E���(��R��QV("*�,Q1U�@DYX�EE"��u�w ���*�TQQVF,T���"����(�(��q����#�}H.|م �b(H���������6��9V�O`s���^�:{ú��s�j�uX�y�W�<�" !����3������$����(��QmL���Q,jP��@�B�=O���y2{�˿}��-��/�⻹�q��O/���}7,���	B1?o�ƌ*��U��/����r�"���_��t���lsQ�$D uN=��(�������%���a�t>xi��]똔|��G��0y�9��k��N�ku�� /FD��(�������L�����q�q��uI|���R�R�D'�{�n���R|+d��"$`�(��v�N��{���N��?$�.��F.|^�̸ZyHV�*M������iS.������b$���5�F�^�x�/��|�0���Y 	�'���EH�Z���"��
��[-� �w�'to�Hu�5	e��j�Z�
j��H�jS��������n��:b(�b)���aDĦ��0����a�� X�Dt:{�1�;�ds�]MI��G:9�BV���D���FX��C�*F�W��,
�
���dRa $��Z��5����9�<��� !�bP���P���+�	ظw��9w��g���Q{�ل�hd�0P�EU Ā��� �(!x� ��lJ��ũ��W�Յ�b`e�X��B�M  4?	��i�:���كb�	]f����X�^"x�|�H�5�! �|:L����W�{�;; � �LL$\L����!�ɟ>r�s>s^ibg�f�a��dӦ�t��Sf��R6�e����u�`89`�0/p��jj�d��AD@�%�Ck�&��wYb@=�u��d0�|֢Cs����/�y��swOC���x��g��<�E�S���	���H�,J�E���q�۫up �\
�D��nȷEb���$����#�݋���t��˒�CC�c���<G|E�f-�.� ��6|�(�n�JI�@����t�ZEM�%@��I|k�VQ0�Db+���y�h9����i�}M���waS�_��z~c��h̵P�v<�Q3��i��Ӿ�Hs���̒� �y{�H�����ۦ8%��0�� d�d@P��Y����Dp��p0�u���ל_b�W�z@xO ���������ޟ#��]~z��~͍�"���XD�%@��]��8������*������;1���xJ0=��A��[��C��?�޹��NPP�['C	HeA�,��~A�g�4��'��y�̀s��Z[}ą�̪[1ǜ�kW�G��ir麞�
��+?J�q�q�c�c��KU"9Y��0��2.�!`ʭ L54l��͍�k>��!�NV��X�}f!�y����z�4ܒ=Q�\��]wax8E�w�o	�H��(2Or�$h��P D���h��0�d@����?�\N)"�T��Z
C=e`A��K���Î{�)�p�v�:��q9����w�Ȑ��T(ȃ��7 2�3D:^��y `�8��h��M�+w���a̔5��".B� l���cvu���eu�雔�U���~�����o��!�@�@1�z�g]��J��gɚ�|�Eւ6��i^�� �"�@��hj$"��
S��Pf���je��$�|6�{�G���^?
i���kZ��PI��8�Z�f9�	0�Yd_+���~'2-M{4i�٩��$"��>6O������<)�����>�9��w;XpS���k�rbT
�H" t���#���O;��ķ4�S����a�@��BG-���5��"_:NF.�#�G�<s�z����[W��%��V�J.AX��M�6ۆ�ā$3�a4F��z1l�FE��RIa 6Ғ,(%��E3r�;�����{��_���S�g�}��
��*xAF�WAp�T}ǥ-� POd�$�H��"�UƐHO�s���ՐVL�3!��<]}���"z^^ `�����DX� 4�`�s�$ʜ�V�id��]�&���2�F����i7��|�̦��5��퟇��c<�{Ts&�3��!1�D ����+`�:Q�!E��d�w��&�ȐRwW� �TҊ��G\�
>��H�L(�p2yc����{@|$t>`�	L�f,#m62����P~�Q�H�ªH�,C� Xuɐ`���>���q���,�{��s�������o[�Z4���E^wx�_��p���4%P�zg�kk��}FsDBD8�T�F]e�R(j��;_��F�p��8� �"Mk�lmƜ�{x�v]+E�1R��2ӽ8rN
4`� !h[5��ֲe]c�E_���y�~W-E�7�ޫ�x3��B��a*;Y�-�~ߤ��ć�d%�e$F�s�U0� �!�v�P��-_��Ng���A�P4���h��lb�>}��T����/9��22��n9^N�PV'Zhx�͎���|� �.t���
CE4�,J�W�CI�2�(���Y�[-i,�,��b{a�y�������q��_%�y>pU�ҭ���kt���%4���1A� Ex3�N
�2^}���yC��C����(�H������T�- dUT�"���e)MB �¿rp{�Y���,���g��7�cs������/?�>|%�����D��5x����B@����Y� T���`V!]��Y�P�O���IՌ�����Y��՗�&��'��d(<�����.EqD� v�D&FB�$$)Ji+����O�X���k������vJ�K'�~�;����e�|4ۗ���3 ��L��ٱ^�r��! ���j��]�i�Eƨ$���x Iu	⨲��(Ӏ�ڼb�g�HhP{�v�p����� ڀ� '���3��U���_S�k���U������	y���ň;�1"E�|!�W0)y�
,-�l���v�M0���M�|��ȹ�y��6�a�%����B,��5�I���r��8��&��C������l̟|Å��x��|C��	`�XJ���e���)�͘��3�6#�8������s�l��
�3�?s�����-ajE1q$Z��4V@�1C
 ���Ok!�L����z����[�#=���,��u�m����x����~��7�z=9��s؀S�
"�A;8 �"B`�dT��Z�j�o/����%��[
�'/�����;��|��
xTz�� ���(�`�8X�_9[�^� ��N����Wl��ʾ!�y�����,fD	b�G�>`X@� �D�"j��KARVD���8 O���k��'Ʋm��>��|��h���ί"%{�)A�)ApK'9����疚�����M��o���;�����"=�^3��ɀ6�n*@*�@����Y"�{��*��E�"w�Њ(���M$�G��oE[락�)�`L2��q��Pm��L�� k��j����\��$z`��_�Qy�~�fAiu�f�	�$;� ��	�,�����UO)=��T1Pd��a'}�Q��A��[/`'�Y?;��J��U!�A����OO����n��-V��P��I ���N�=��`�lL���(G�XG!E	
��S/���߅�P�����߽�{A��fʑ�����r: Ul�-#��[	͛�t��`��|K!1|(�(y�P���(H0�u^�7��F��{�ކ}��w<��y�s�����o}���"/M		�R$;���Տ������8�'4-E�*�l(��x#,X�	%b�(N��'��� �|z:�9r��,W#��t�f��i�����#��^	��N�zl���^~��_Y�͹�+~�p������ �:
�"�l��t\�j"A$E�!,P�AHE�����!��ȇ�+�l g�:�_��[��������-����U+��w��J��(C7����jX�Db0����z���3�Nk���^^od���a���w��$S����.g�6F���v���:��8���w��ʮ�PM�{����BlʮLR�(u��`��F�$��=����"+?��n��F�$8:�an��`YIt����(���V�
�C�P���0�0֏��շ��������L��*M�鸂c9�3{����Nc���U ���20Q���y��(!5)� �B�F���[!HKbRi[�=o1�e����]��A 0w���X���P�Dl��=�7�MiG�=ϰ���ެ����' =���fx� FD �!IQ.D)��UI���P)l᪇�`�OGW�g�9���=I���CH�E\�1@��	�j		 �^.Ӗ��o_��~��v�'��:H��������18pH1�#5JZ�D]q#fQ��%�gb���<�JW�g@Ǌ�_���D�3��Śk�|%��(9K��#��@8���X�,�`9�)�v��p��lF��)b(�"�����$!���&�MhR!)���$a�<���N}��|��q���:�;�;nb���w����,�L��G��X�H�"��u�����Y&�`��F�@��-�'�@j pR'�߆[�'e��(f�  �K"%�@P�p���@��ۻ ���<�c�02�^��Oq6pǟ�՗��T ߑ>D��"�I"���T-`r�OC�s��W��Q�� |9c�ޕ����_M�:2a:S��7��/�`h��n.Ο������P�&5A�L+�dpHj�Y �@�dR�F�ZŪ2w�;�	�#��|�bfS�}x3����2lO�;/mshzY�%����/�I�@bt�`�:��:�4d-��VN��r�I��_�k`���^wz!=�?��XuA�$eG]��,X�
�R��덽������7����EW���df�Sc�݌��"�'d������E�P5b��c'A�Y<F9�60�J#=��(���Jș)�yޢ���� �|J�z�
�@��=�9�d@c����9��OE뻼�oT�H^>5�L>7��ٿkO2�; �Y@�9�[a�4��Ȓt��E7�T�_�;?۷�G1i��k���������9m�4��5�e�9ik;�(HA��B�Q!8�Z��4�V`��*~M�3�/��w`��cܞ���[���^-�;���i�,Wu��"0?z�@�=�X��;��=���T�ДTJׁk]N���=ځ��X� ���7�Ɇ�y�o.3c�{�[�7p9�;Y`�"D���[+>��$�������1���������*)��n���#l�_�����s��_����#��~�\�Jn`����A�"���0/@?bPw1 VAE��0@��"}��*�Q��rz|FRX/�z�a+ހ�����t>`�Yf�>�t�8�c��װi�3bϻY}Q�FLX%e�����ڿ�n9vg�y碖9d�(�� }��u�&������M��t>��yՕ4kA0R� ���f���y=�}dR~u��X,M�:��`������?efA��|[�_���`GLq-�4����T�Fo{K��\���a�����o3�Ci����dŸͨX�k}6��Z��ԀB%��`憤�Z`îP�xj}�҄ZTN��8��
��P�қ��&e5,�y{�l�<:E׿{�޻����n
�k�}*)לz_k��2�6��
L� ��m�C��P��DS�X��a4�g�d.S�K��h��2��3!36��4ά�ft̕�L�0u���O6\��Vgo�|����������+:��f��9O|<�^w��ӿ<�h;;+��|�H˨���_ü�e��g�����B*�t��@�<!M-�V���V���k5�R�P�t&��b&� ��ͥ6�i9��ǃB���	����[C���ǡ�W�b�x^^Y�Y�5�G�`t��Qq�x7�uI4v^�%0�@�۟���T�S��������w�����9y�%����F1��0I6>;�(F�PL�Ș�b�� �Έ� Ms��[��������)w� Fg|ed��'� V�U�G�n����,�	J}+Z�@�5>܉{)B���X��/�kьcg�+��_�B�	�l�'�����A��̈��Fo8�bl�*TF!x��*�@����X�a��T�o3��Gb�9ͫr|Łz�K�9QR�"'V����A�� ��H p��G����a��7a � <��2�*A�u
��KQa�����	��� �"S�>�	ވ�,T��s� ��(Y@�(@�Edw�YX�օ9�W�������C򑹖�~J@)�i�����|����8�$6H�Q`<����)�Fh|���8�/��7t`i��Ď���t��"���E��1d����"b1�`��\�+�����.�<f���Y�kB�q"H���fo����gK�$dL���:�� ��QM�E��4\�iq���7ν������gM�D��k�+"�>;]X�;�y��1�H���@H��д�IH2�PE�9�����[d�|G���<q��ܬ[�l_���_�������g��G�8Z(J�B�?f�Vd�x��f , J�q�(Z��aa��,�	�/�ƅ�~�("[@s��`���T�P,ؠ��u܀6�8Z�y�kOb<Mjͭ���*=@ _�<�����Ԫ��D!��I���醑p?���t̀[�pP5E@P��R�ʥΑ@���z�x:�� hn�JN0�#��"9OuL ��퀞-#�� ew*aҘk
�f� �%��:S�Wp6������[x����f�@mT�EP �LC>����a���	�P0�k^o�� ��D���(��� #tJS�	��Sr�ݡ�c��(�@i�e5A����(k<Ʋp����Z�� y@Dn�f@� `��
M j��&�,v]+�"�4��2�^�g(�3
9�b���o��R��t��P5i ���#�,u�#���>���:�xHM�	���(�%f�-�"?���-��R	�P9�S� ��D�T�����8��&����D� ��K�q�P��ϠC0�~�y�����=C������*x���$H$�Ă	 #w�PB���E�£A{�$����|:4��� �x�� ��&��� ,!�d! B6Q�� l�;�!����nH>7pl3%��@2A�Tb�P")��WCn�� ��. @�s�%'I���n"6+�H��(�0ӏ�OJ�� t�K]�ӣ ��� �I|fCO�j�(Ą,�&b�\��s��@9Y2$3-`b	��r�(ɗ�W,�2���(����w�a���Db�'T��7����  3(�c'�k���ۋa�5�����;
.<~���<Tp��j�1�ٝȡ�bA�wʬ��<"�TI'Y�7�,�/^S��h��20�	�4��lTӱ���H�( t^� :����� �pj  �t�b��t�, 	$BDSaQ(^
m�����R�� �� @ $@�UdId�B���
��.(sd	Mw)�SU�
�@GH^�(<E\P0pBU���|;�� (����nH@`�VP6C���\��V� p��@��C0�@:C�(�`�y��
ӣ�`F#�5�v9)�5@,��+N4h̪hR �&� ���ʠv�[�"�p��:
�#{�y���l��XC1Iuq��Qj*��Ȇ!��� �d�j;
�.�-�"fM��M�ح�Cy D΀��H r���!4)�e�7��=���6@{��j�\�B5���,m [���k��>\=�&�i�F��������=�Q�]�	A3�Kd�� w�UK��)��J噶H�${R��"2
�H[�B��V�_s��?w-X%P�w��N�lSj��b��I�z�9����e�J+��d���Ve�?o�����G��7[�Y=_X�-��,�{�0 x�<\��j��@���s`m�"���Jc×"�j�t��î���[���-��v(AP"�	[CT����_�ߐ�U��wʰ׺���I@Pb �`�`� �h�'����#!!�A�w��1X� ҁIb!*�X�LH[!@�B��Y<V'ij��W�2P6�i O�P"��n�� �������l�� ���N�Q�74UM��H�Ew_����Y%i����N�<f<I�����"m(S��k�3hB���[K�)O��.LohB ةAV3rP��`F� ��P�n�����H�4�4Ab��H@��Ou�l�b�Q��Y
@�_O��� ��f�C�(&�@֠Di@� <��`Du/�.!Ϩ���5�|A.�@�^��tjř�1�$��EE�*�'� �@3&�"�!	"y���xa�8�l
��q^��̏l\Cdk�`4�\ Mp8@-xc(
�@���<��(@"\�ew� <A����	�~s�6�y�}	�p/�]@�&�euҧ�d�7U�����Oa������������|6s�L�s�T�*�堁N�r���z#h�
�D�>N?��h���E"�RA�*�F���C^O��S�}�n���#�@u{z	�� �D@��`����X=��[^Oa�I�=����õ'��(�Ɍ�;���$�&��"��R�� v�������(a �~��P:�H�(I�P����~	f�g�JT��� R �h(�"�aLfH� ,�6iW��y �)׊C��q�;E <Z��p K �,�.�W�貁��v
�e��luA16�8��FK�m���o0���K�}}�`|�8����~��O�CMd��ƅ�(lׄ����pv��������l@I`�-��*�>�_Q�i02���"zXx��PV��P( 9b��EN�W��˄B���i �{��qP9	��8e!�t@��Dv�6ာA��X�*j�>�û�q "^	��N_��� TT-S��tZ� �~��Q���s	������W�c���1"!UD�2,�T��Гhy@�	�2B��d�[EDY۴�M�_��u�@<�;��X"���`����_�P'`+��ȬD�%���� � �D\ ���
�s'2�0�C s�T�g�r���;=:v�8F�'��T{ԇ��)D�V1{��`b�F����*�@g�l�D� �h�\���d�V�8P� �b Y �(o
��$˅K*+��f6@)�ct�y�� �t�Hl!��[�$V��@K�j]� @D�� @,1[�:L�t.d���,�ZȀ^� ����@��e ���en��M\0 `.���a��*,Q[��^�"#;,Z�?���kr�dE�����17�x4��n#$�����2��+F`�8�!ɉ"��E���倦H��c �UF�*(1Ty�d�<\�Al%��r�2��#��vpz�p�ӛ�I�D3�?����T@������KO�O�sv�@��R���5T��XP�i�*��`��@"0�I�M����m�s ����C�*��([Gp������u�Bú�@2m��D�������������zoa���"�ϫ��gq$�~"N�	VAXAU�bB,"0Dв��d�"J����(Қ\qR�b!Hv6�0܅	�L��[llF�&o����ƾ[�.[MB���B��k �T	�@#K܊� P�h�3ryT� ��M_����pOq�ri�k  ��el&� � 	]m��F�-�����2�c��OP�*�����K�����GA����3+� b�rg�j
D$�����j H�����|om�l�����i/����z��g��.og��'��/�!��h��/W
�*Q���(2�,X���$"@V(��ĉ�%�{�g $�i�y�#��:��->�-�\�x�:�( �S$&)�n�@��� P�
B��]fԠ^�U �� x " m �W:�oY� �43��A֊�`E�[EZU�
 :�A�ʺn�$�WI�`"@D6 q[�����@��!F#Q�d]����+�T��q�EU���`a�^dQ6(V�Y
x`<�$�/,����!e`U�)u���'?7NwQ�S�2��HI!Bwa:�6�Iw�ܠ�;��ن�fr00G~$�Ȩ�u��'�CA��@4���
��J��t�7.��UJA�9��I	�!$t@P���^@I�n@2 � �J �P6͔5.����B(� v�P�c5 t�CR6��r� �p��$���u� �<��8�O�������eykq�`�O�m��HI����B�@�aQV��ƒVj�"�E*�?M�0 ?��,��e�O԰���9�5Q���ʔn�f��r/ DI$|(�f99"qW5'6�� D #Վ��� ���P3E.p�\�9)�M�\)dT�4����:?�"h� 1&d�YU/\0B	a��3�H�P2>iQ@�\����@0�A�� D�UT/��6�~t��7^����eM��PꣷGb) ����K�HF(t�J# ̡�7V~.��C��ְ�"#,c��W�u@��;�jP ���	��P@W���OJ� �.� ��� �* ��h�P:p ���G��sME0j(_ �7r�g�N�H��!����A��UL5�M`D��E0wR.@��*��~U����ó�TE��Z�d�<F�x���Fp@�CҰ���IQcH�UPb���h�`Y<L̴��d`�H�>_��p�R, �@�� �S�Or��et�.y�����}�j�p�|D���[���a`Dn�%Q�$X@� �%��P>Ү#��9Y�ާ/�v�0xv��r\��yK��!��5	�˙΋t������{��b�9`��B�ģ�������B�U �4ȐU"F�P���PdP�@R0�v�*ԝ��R��J������/��Ú�7�s/�c���q+���/3��0��V�D��H, *+k@Z�(��d`Z�$Y'Ъ� �)�8H
d�AK)bP��I��lA�8�#@���°P�+V9-��&	��/��+��=F�~+���O�݈�Ǽ��9��#���vB$��E 6�;�(b!�o��,��Qћ����ZRr�"��ǐ�� . �PHe�C����y���{,��������w@xuy嚄FdEQ@@1�IO6d@ ��2"c�Pi�V*��H;�L�ϟrj��e����K��`���4�Y��� c��B�b
	Q`� HH)2F
�F�ňT��)PYJh��������ʱQN� r���o�ǫ���*�K�>f�Ұ�̟E�;l�!���U:�`y�&����2�/��P�L����a <�,R0�Yx�.�2bU���V�మ(PS�
�mS���@P��呥l# VH�B�_�ʬ$6��Hz�d��*��^��~ ���7������a�b=����+䢶렮�b�(I �;���US�9�Q����,���"-��H�x�2��(�>U������y���E)UJW�nzW�}���y��:���ohhAN���L`b;l�"���.���+	�R�`�*�B���8�K	��
���=}<�/2�~��)`*��$�AϯUu�Qe����7&��%G,?3��'���M�Q(!��,f���j�`��!�!��\d�֯)��}��k��$�"xH�~G��zb+ߐ���9�d:�Q�j�G+��YT�	�TeU�?���-�
�I/{�/�sm��n�殣�aهV�QE,X�bŋ�P�^*L��Y��	cJ���~�k����`���c2V�Ç��@θ�T����w
��2o�/�����:�)��EeJ����A� h5Z1R�?�� ,�
�~NWHє��G�zo��?��n�]�g���w�`�&�̷R�	�ˉ
$�尲��I� �DZWIV��}���=�(�?�E��z�"�	���zP��%%��H�����߃�=FC�۝t�Q|d;_�O��U1>�jIh �T%B��$�@�wd&�C�倵)C�m�l�㥣��Rq)�&r	�"�&���I�z���_'��}⁜�x	 :����U��hA��E �0$�(c����8���m��M�y�ٵ��}�������:��חMBN�rZ�#��*�D�U�Y��P����m�*���'ek-��i�v�	��`��۸q��L<�l�HEQ			>��`�ˇ���-�L�p�S�dxd�:�_ĭ'�͏�a�2��e ( �Nr��V ��|��h�@Q�qNa�VR�,AK|jr���Ao�����s��hȫ���C�C<��h_ P"���F�F� 6_�S�}aZ��+�����޲��CŀQ�v��[�X�H��ve�.��)�vF�WZR&�H��UE���A�M�>������@�)�{z�O���E}���m���s}/������x�;N��y��
�.a@?�x}T~T
����.�%���������V�b��������yO�W��L�e�_���9w~g�ɗ����Ƕ���������Ȼ�H�7�h�X*ATx),$�d��0�b�I�,	A
�P^"[��W��=���_��-����(�RǇ������t(W<=3c$ B�`E�Y,�m<�W�{��q�I �I!	��O�/�}��;�yA1��C/?�����;�z����<�^�&Ҽ��WU[EB"2��Q�.7�_5^��'�]� �"2���i�}�0KCX�o#�����^X�:n�m�Z�������Hl�)-aB����	V!B�wAw6��������d�}Ɵ��v^2{=���?à�?{���3�����B$�QD�R��|�KYJD$��{���9s���]w�v?8��v��7?�X�*�+-g�~�O��-�tΙ�:ۇ����ñ�tD?Rs�Ղ)ZU��\�H"�>́��Ha��;�qX�|ꪳ绍S�Z�M��+Y�`+�0D��"v�:I�A<�G�f̐� �� � 0�!S�R���23�.��owN�3:\�*���r@�����z#��*ԛEB}�u,�+�s~qb����lC�Xn����^��1�{��翢�0.�����v��b
l@I��E"ZhaPH�@A�=�I�mRDQ�K@�fjӰ�9��Zd�<k�&�����DN�+��v������~�z����o�ߩ"!�8�,�� 6���*H,!E p���^N&&Nz�Yz^&�S֩�bE�P����"���/�)�Yć<x���Pq.���l4�'U���=A�I��(B�D�dL ް��*d`��Ƒ��!K�5@��*���`0�N������	��k�{Tj+�`Hz�(�pR�x��(������?������X�Iqd���	�1�L�����?�9?K���7��������5i އO�Qʽa�Y���>��_!�e�!ݰ�0xe�E4O9�Vq~�������������=V�؁�^`*4�	N�Z�P^�HD���������>���g��S̓��zwu��2��(������9<$���S?��J�"�` f�QB <�PӿY����s};~O������e�a�X.>O�s_B��[�o���2���bA�9�{�"*-�hH�>��a�_���
n��AŮ�~H\D�&�i$q	��UE�9
hxd6
�5[�5��^��K�d` ����o��';�����7RtfBd)	XD}S폶��r��, ��2�f�-��.�+s?���_�퍍�?�00��KT2�E!D_�;ؐ����L!�?K����~G�u2���>��������"us��P�!E����������xLմ{f����/O�rr�toRSf��MI����X� �)%� �����C25^��1 r~W��9��f�8ҭ�D3�X	��(Z+/ �6"��'������Yq���!:��H
���Ü�P�E�#�2���������|�k�u���x����y�T�暂,!$�v�1� ��0��D�-k����G�/�>Zc�3�W��^{�!�D:���h���w,,�O|�����|, ��o~���MU��H������澖m���o|xq�'m0.� @!h��s�md*~D׻!�}�g���,x�z??������z���M+��7�8"`m@%Ed � ȅ�/�|2���>>�N����k�@��
�;vGgd慔}L��i���O�� "	I��DQ��������ܘ{�z ���HH'}�=e�:{�o/-?W�k��:��B������Y�^��oXc�Ί�	 ]��������g���.�:y�T�B�H�	�Z�>[�������v
�9� ���\���݆���K��F؈���ٍ�`DH����G����^�V|{������Xx̵l=[��wݯ'|x�f��#����!t�B����`a�����;8HX��
n�`���~
`z�뗤��o��z�~���#kz!=,]H,��uĉ�e�R!�y�e� �Z)Y�����/��������t[���vnv'���'���?�gԡ��4�+'�����;�j����?�6��]_h�"!���`,�;[�=�� J�K0	��`��Ռ. �4%��C����b���'�D_{�oEn6>���Wc��Yu���������vl	l��E��`0@π�Yd�3+���U�^�8�5�[�~���n�&�$E����_��r� ���Nf�{@@�=����ҁ{@�����J(C�x2����8n%%4T[� �>~����>VT�����GXv�'���o{_��co�{8܎���hD�k!��ZH�<��LA

)
�(Z�)yx�'ږ�_�[��z+��'��f�lr�a����/bv�j���F�3��'�~/�=���/u�Ti��gb�|�����J!�0�H�D�����N_G�|�O��/�������������S�����&�7�J
B'8݅��/�"b��Ci�W:��{�K�M�_���)������6�D���/��BBD8Ѣ�'�\/H�Cqb����{���zV�L����.������ro�v�f��)}�CǷ~Y�y#MO��w�Jq-bL3R��$$p���s�����K�%2"B `���v�dz�&���E�"��+ʂ��x|�=��v}�FN�ݴ�C@�� 8�I�B AA��@�2pHn��Ʌ�����nBo�8�#�~]�}�i�#��@p�--���!aBW���5�#�'�����Z���M�R����P��O��B�Gd ���U��ͨK�L�<�����(���z~������z��-(��PM�����AZ�)�Z�����>g���_?����w;/Q�� �4Ic�<�r	���J�.��,�) m������}#�N���K{^��A��j�IbF�dN�Q -�4-D�:"2�����s&�������R|��뇧�A�zO��?���������m�A�Y��*� =uH�6��2�9��֣�zj1��� �k�5!���5P ��:���{�IȊ�������<e�w�)�������u��kAc;�W��!�,�����tc����cI�V�@���ϋ}�py�9��0Iq2�B
�� �	.Gݢ���\��_.ȸޢ�r4�0  d��ă�������B����z�~$�ɜ�x�~�{�ϸt=��c#�0;�A��K\�2�]�Ah�!�E*�"�v�ˁ�� o���ޭ�3Ҋ��Qo<�S��wq��݅!�����,>9�������jN{�=2 A��
?��7�A����J�=������q̖��RX��� ;,n��ZP�V�@�>�$Az<���~N���f�o@�j
l��aa)d�=k)#u���ן��p&Y��Q^� �������1������Ϝ����1帼Tw�I�ˈޝ�Źp�q¨U¤DK@P��?j�����`SE���g����������鍩M�B�e6���F�~<�� s�C�{�������0}��������տ���?�w[!���ٶF�$߇�٦�JB*e�Ep��0*~�-e:n�&�e"���8Pl��d�P�AU$�=OW�����������z���@�p&C�C�����cN��=��#��)�L��������ݺ��5�W�?}�k[����}��X��>VIq���iO�h�tP��iPRg��
�oj���ַ>��M}���-����7e�L]c�6<�;����=s�5�q��@�D[O�d�� ����O�g��=�\��_gz�'9�)��F�	n�w�/ �B"�"��C	�h�
 P����ð�D=��s]��*�p�e��D��XaD��Mx�=��(��OUl�޳��'�qwA���F�e�>�_+��ﷹ�� 
bB1��1h���@뢵t�� �1G��m!{�@ob],�ԁ�V{��|l�!��s���Ƣ=���#HԤ�4?�kv�?���}�NW��>�{��r��L���P� �MkX 6yߔ\�a�}M|�>�x���������(ւ}�L�^[�p�&q k)k ��Z�!P�$�A�(	K��-�^��eqE��r��c���}���rم��(�I=C�3��� bP0�(	<�|4�?Qe�l*o��va��V�w������yo7���P��BB�@�
�V �ʨI��s�mc���}(�X�q��
�H�PJ�=풂�(*���1��k,X�((�"(@D#"��,UEA"(
E+�"ĲU��J�֔F(���j2,�Fն*���D�~e1��@��|�M=�_X$ �wyu���F��/�V7H_��^&��7V�b�.5�9�jܮ7�[7ԇuƣ���]s�g;�}��k�X0�+���,�Z��+X(p��W���R�L=����Ԕ0��H0�$�'[6������{B������%�R���p�ΰvU;s�,*�{­^.��sx
���P����s\��V�"b?�c�a�t��K��5j�@��{�P�6�w7K�4�1��^7 H��JA�	M?Δʻk�l0L���̒��U�Kn�K�\�D���GbP�����"@�W+�!j_�<�������t4uqn��Z�4�5�(O�+��"�W�*��C�"�H�� ����3584R�2�L+*�?�"���\�uԈ<��
���ވ�5�Ș�)'�g�òph흸J�t���V!f/�NŇ�������&�@��P܈Ƞ�i����ҟ�[��Z�T������O���(3C_�e��BƄ��%����8��<)��s������y�_���K}Ir���Ql3TFH�W��<��@�s��G�1���U���z<M\�+�0��Ֆ1��S�8�#�?����J��E�� ([ho�X������~���מa�p�sk�w�2P(zcj���!"zD9�0p�[ya;c'鏀3��qI?ఋ��'���?t�TH4�33fiՉb
,+(RJ���OBS����߫��uӞ��53��ך�S���`TV�	G��Tl4�Qm YJJ�S��,�_���3�ai��&�8�1����٭���Ս�����W������Y_Yy	@��m�� � a��`�%t����%Є����o�X����7u߿�E��0E����/���k<=>���{# �   ITr�Jl���_O��)>$�����Ϲ�n�2ù�?�K�,��2�X�@��$��2u�����])����j%��)�4]C�TȈ,MS"H���bD���-�d*T��b�]|�>��̀��e&]Gb�
�7 ��VD?� ���T>p�^2Z
*�����<�p#B+O}qB�Y
e''P�m�0��m��iX��|ӱk�����<Må����f5$w~��Oop�31HDh�(B� �����w�VC���V�����x?W���q��[���z6���Bz�2!H� B��
�VW��|�������|�*EX��wjs(h�g������;?���������B�7av) ����?�i����,�A�HT-��S�N�8C�b���F\߉��ϗ��l���mw������|��9GK����0��,ĂA<u�@��T^,_�"rx�ԛ������8���ʺ��/-�P�y������Sl�̣Rc(�H�;�M������Ǯ/�_����p�����y�u��߶���v��ȄYU�J^�5�[�:��5i��O6#c�|�_{��;��"+�dr����#��C�]��f�|�7���~��rO����zM%"���a��(�4����J20A�H����f�s�8]�%�w�7��=9X]��RxO��'�w�l���Z�EC]/����T�YX�"� ��Cٙ��S�����'yA����K�R~f�u����k��3!�F�����B}�,K5+÷�>�����k�.u]�#p��'���<����?������w��ĭb�5F J`��(��	��_�#�Ƥ~���FO���-��(<4z_��/����K�����5Y�f,B��2͉����=N���{\~�׋�[�jQ1b�	����B�e��$a��(d�ݸE�C�4b��E �l�p�����e��XRV��ݶ�5 � �@<��XA�<׉�a������C��zm���TZY �z��c$PVM5P+�O�qu�'���w�¼׬��������_���;���W��T El`tp{���K���?�YveC>U����,�z��ۑǤ��i^�TdB�/-�S³fu��	I')�%���R�1��z;�����*��j�~B�u�&�W���y����9x��P����]��+-�~�oW�z�l>v��^�W���?���D�0p�{ �@
Y(�(�,Y,A}<��9��u�_/����?V:��|��	�~����� _���������T E�t���`����<�n��O�Ȫ��p��O�isj�/u\˗y�0j��h�eJ�}��	�r��-���ID�  D�Xȥ�\ �`�@k!aC�>$֍0A���PH��RR  �,���=�������r�r�]3>.F��O�ɑ�p������y�?;$vgoN��z����C��ڔ�}p a�a�O��B��Fo�����-����p9{�N%s��9&���[�M�7�)"ŵ��!�0@ ��4�� ��{���r8��b��a�Q,����3����]���T��?ٿoe���o:��QCw�w���Q:��l!�[Y�P�0�>X�����m�[��Bt��1����0�!ؐ@�`�9�ˎ��.�?^��LE�h�u�#MgO9|6�>]��wg��'wj��|�J��]�X�����?�G���^����#�j~����?'���������S�{�E��=x࣫ ��
��'Íz�~��V ʕ&~����z�����<���6����e���t�+2�/��}Ƹ�����3)�Ē�g��fꕅB��\�T9,KA$&U�����d!x�0�녺��aޗ� u&����<�����$ti�T�'���=����#�R�I��|��k:<����ҿ����'�C������v�
���NRVn��.�&�7�`���fX�p?&vpq%�i�@�	#ff�ł�FXJ �0�AG}4���T]/��U���������KZ��gciW���d��E�V�h�K�t7Ej!����R�+52�c�U:��F��C̶����b�7:����uF㮢)i�G��[��%���IW����`a�
#�ſ�>/�@���߹*�;-��� ������88$|V���y�v�|��W�H㺲l����a����7�?&��m��:���(D����L�D~h���P!`!������i�̋!��02!bP�	$���۱ӎ~ôOR�ʆ=\�U����F�{Hx�!���,׎B�"g��^��iJ�������9���-Q�L�*;I)�i_����·����FjGe^�K5�� bJ���If�4L*�ە�D��i�wb���5h9�P~�������Q��@ِ�T ��Q�Zȯ���n��m{h�������5A���Z�/����!�!@ �Q@*Hġ�(H�N��yy��������Mp��,lA����<�3dq�ʁ��~��[�MKۡ�9^h��H9�sl�f��̂��s3f|�uM[}Ve���ֲ��~�0ȼ�F�̡U4WR�&��\ڂ�������lkL:��|�!`�?.v���1)@�B��V��9�MF6CWx�Y�R:�놞��w��O��4��;s��N
W�� Z0l��4��@ ��O;/39(��}��㚒��c�HY�hgV�t.�?Ϯ9�|��{.�j�f��cڱ��i�7h��d�E���^�y�R�]S�N&i]iZ�α����k���5h%�˟�b����\޼�O��u��
������j��J���6������2�A�]�Sk�y� �3��jV/wt��д�b����������Z�Ǔ���r!h��ό����r��t�_�����=7��{,>�Ap�
�P  �F�*B�>�(Z
�!"�H��A
z����ݑ'G�����n�ʱ��J#���uhn��-t`��I���u�m1Nk�R��[����Nȴ�V-^�"�?ײ�Sɡ�f���.��s۱��ȡA=Z[�������O�M���\Z�����^�Y�}��#t�t�a��V�x�M��z+�sX�o�1.p�J.11�X%m�8\J��rI��ed��"�?�k�9��1� s �]�
�o�E����ܹ�ڬu[����޻;��(��:A�~���O����<�َ+Se��~�O��}���9SBX2X  O?��ЄA5(�#
3�HRA���� �=@P�"D l���ᇈ���)��US�rk�I�W�SSH�����~�N״�=����Љb�.y���:�웳��圊��s��p�/��^�%c���2�g,Jvd�*R�4���aw,�֫/4h�iʋW ��9��Ky\��rDњ�M2�B��3ep�٩�ܘ`i�Q]��7�e{��l��L�����,�Ϭ��V�ۙ2���4�LM�DB�c�~rZrȈ��@�2-�Z�T�i5�����g�i6���,�jjO�k������q�kO6o��aY)Ʊ�wnz����顰3���������	\*B�]��Dp�:�c��.�S�'?���WI��'K�H�Yԛ�~�f:����9d���M�^�5���&��j�6z���VX���y��}j�+ɓ�pVE�o�5�i�+���,Ԓ��Mf��ӱe�Tj�����ӉkO�`��B�Cy+�Ù�UoN���t�������V	[���,mm�B�T�蹪����`~��<bȟ5s���{Xi�=-צ�,���Gq��z���!�5��F�xa���ˡ���<�>P t z�"�gQ��5l��ꑑf�����7��o�9M�����U�{��Eu�o���Od	Q��(����3���ٌk
��I�?������Ş7�o�ORr�n�*)��@��I���=���}J��b����#$��f�5ގ�yX|hv��W�,6U(�T����{�9�-o7�}O�����з�1,cp��7�5��ҥ��ͪꦍ�%�����r9l��z�nw��^z:�{:����;J��ug�s��-ZX��k��E)�L�l��ǐ�Cez�U�si�����8����+D��v{o���K ��ʘ�f֧4h�n]{SE=�cn㢻W1E%�/*���f��}3�{5^��}3��b)�M��e5[�[��(a�j´�i���no�9t�?3Ӆ�r'w1�8~��E>�|���;>���U�:���~*;j��y1&��������-@��5H��%f*�ѵ������n�ɵkv���ĉ(0�\����א^�F,���������ک�H�^�S��[�6�����w`�࣡�@� A��;�0��yww�1���d�]˙��RnHzS���z���.%���4 F�@]L������sn��W�O/9����lsQ�u��{���"�v/�9�S�͡�gܔ_�Z�����?nO���?����79X����~~�x ��	��^�'��<�Z�zo���9�/�i8���[ƫG�z�oc�ȼU��xX8/���F���3�KHp�F.���Z�h�Ev�+z�8ַE��x8�J(��p��y���(�z���&W����u��Zc���']"0q�#���@�_z_�$�0P>M.�RTI4��"� H ��(��*�"�*� 2*�"���A`V,
�"�Ha*@���H�VQV�e��PU ���I$""3�B�QRI#"I$PQP�@QD�P$PP�YY$YB@@E� ��  @p�e�4�1T0R`�b1Q"�F)/��_G���Ϋ���ڽ_��_Ku��O�ۛ�TDz	;ddb�`��"��b�Q0EE��4�t��X�`W]�QI @��p��.�.�J���9�����Z��}�e�|u��}�gGZ>3��+ị:Qq�۰{�;9?�oA\��^������|��p=��ű�'��v�1k[^��h�Φ�U�������t�\ٯ�Vm�}fo`��Z����NydMZ�rw��/�q�Ik<ט�;�ˣN�O�c�Z�f���V��Ӹ�ͼ��N�����c�z7.]��V.���7]��`��?�A%��$��r�=�l`��jM3�\�LT� �}[�K��YO��� �����=�T����y���y������Z�J� �(���1���e*)UJWa�b`�@3�d)�E
Q�����Dj��x���UJ^-�R��R�Bf"�8�l"�$ �őL�JPY����{��?B���7�_&�"@@B��
H�(�����"  Y G�D*(��*aT���&��R��A^v��W��.v�*D@$,������D��y`i��݆u��-/�n�W#���e�����"ɁIu�]aj�n�'K~�^�gva�'��;���AT��/2^�g��c��a����Z�f��������ד��%��G�u�c{zP��/U�;_�|����(�%��Ϧ�FЀ!�{MO-7o�r��"���n-2�6�q#W���8�$���͵�����I�r����-���%i䴉�0�� <��!4�J���4�l��.��A
4d(�G���7�3���57�P
�F�~EU��!Ztɑ	�+>�ZP�lk|��||_�b�9 �8E��^�e��򪁐�<��":�иϡ`��U'�PO�[��<u}��b���z�{�Ғ�������[���y��}��9}*�Z��������	]!��]�0��[XLa�cЗ�G�2�t+���!R��9A�k��3H�o"P����ftȼ�"��"�I���cq԰��U�o�f\�l�`�C/(��$s�^��V���!B[hyR2L~d�O��B��7i�1 �1�;y)�uؑ�.�eA�^�8"Z*�nɌ?�i�~��r�s>��eF�8G��-��ܰ�Nx~��8~H?P�ӌ>+��
���K��M��������]�P�pc���	:�"+Kad����6ͫ2P��?��7�=g�� �l�2����V��y�FPx�����v�e���
r�o��籎x����86p�U !- �g��qz�B�M���(GJ��W���Uǵ?�8�De�F¢@���'����ic 1�z�Br�k�~t��ַ�i�(�)�k�D�}w�|��`��<��]��������S:�T�W}0n'?�|�e�y~|r;����^��7/�������^/*��~�z|��_U�g�f���/����� cS��/��>�!��8[֨@�<��풎��^f;i���vZx�V|5.�ed�m�D+.�e�d����7\m��{�$7�1�G'�p���(�UwT����oؿ�	�AWO���F�j�Y�,�1{P�O�D��s�,����T!*)�f.i���h��eU-S���٬U�=��u�B�§�PYr�����������.��&���g�z�ẖ�->",.�X7�az쯷���P�[L��܇��Q:ԋ6I����Gݥpd/S����=���p��]�:�]�?���:8�\�1Y	bn*.Q����w\�3������Pҋ��[ <{��00*[ګ�������zj�L0�A�"� � f@�n��d�/�J�'�#�ttg!�q�v���v��b�3��Ҿ{n�������{�[��b���{u�;�~.D��|_�����;@��FV@@�����م��lp�������򁠇���Y�e	c�_�-���z�g��H>�NF�pwE8�o�#��Q?�]��BBX�nh